--------------------------------------------------------------------------------
-- Entity: acia6551
-- Date:2018-11-13  
-- Author: gideon     
--
-- Description: This is a simple implementation of the 6551.
--              It does not actually have a serial port, but just behaves like
--              it does.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

use work.io_bus_pkg.all;
use work.slot_bus_pkg.all;

entity acia6551 is
port (
    clock           : in  std_logic;
    reset           : in  std_logic;

    -- C64 side interface
    slot_req        : in  t_slot_req;
    slot_resp       : out t_slot_resp;
    slot_irq        : out std_logic;
        
    -- io interface for local cpu
    io_req          : in  t_io_req;
    io_resp         : out t_io_resp;
    io_irq          : out std_logic );

end entity;

architecture arch of acia6551 is
    constant c_addr_data_register       : unsigned(1 downto 0) := "00";
    constant c_addr_status_register     : unsigned(1 downto 0) := "01"; -- writing causes reset
    constant c_addr_command_register    : unsigned(1 downto 0) := "10";
    constant c_addr_control_register    : unsigned(1 downto 0) := "11";

    signal rx_data          : std_logic_vector(7 downto 0);
    signal status           : std_logic_vector(7 downto 0);
    signal command          : std_logic_vector(7 downto 0);
    signal control          : std_logic_vector(7 downto 0);

    signal tx_data_push : std_logic;
    signal rx_data_pull : std_logic;
    
    alias irq           : std_logic is status(7);
    alias dsr_n         : std_logic is status(6);
    alias dcd_n         : std_logic is status(5);
    alias tx_empty      : std_logic is status(4);
    alias rx_empty      : std_logic is status(3);
    alias overrun_err   : std_logic is status(2);
    alias framing_err   : std_logic is status(1);
    alias parity_err    : std_logic is status(0);

    signal soft_reset       : std_logic;
    signal rx_interrupt     : std_logic;
    signal tx_interrupt     : std_logic;
    signal cts              : std_logic; -- written by sys
    signal rts              : std_logic; -- written by slot (command register)

    signal rx_head, rx_tail : unsigned(7 downto 0);
    signal tx_head, tx_tail : unsigned(7 downto 0);

    signal b_address        : unsigned(9 downto 0);
    signal b_rdata          : std_logic_vector(7 downto 0);
    signal b_wdata          : std_logic_vector(7 downto 0);
    signal b_en, b_we       : std_logic;
begin
    with slot_req.bus_address(1 downto 0) select slot_resp.data <=
        rx_data     when c_addr_data_register,
        status      when c_addr_status_register,
        command     when c_addr_command_register, 
        control     when c_addr_control_register,
        X"FF"       when others;   

    irq       <= (rx_interrupt and command(1)) or (tx_interrupt and command(2) and not command(3));
    slot_irq  <= irq;
    rts       <= command(2) or command(3);
    
    process(clock)
    begin
        if rising_edge(clock) then
            soft_reset <= '0';
            tx_data_push <= '0';
            rx_data_pull <= '0';
            
            b_en <= '0';
            b_we <= '0';
            b_address <= (others => 'X');
            b_wdata <= (others => 'X');

            if tx_data_push = '1' then
                b_address <= tx_head;
                b_wdata <= tx_data;
                b_we <= '1';
                b_en <= '1';
                tx_head <= tx_head + 1; -- TODO: Bounds check
            elsif rx_data_valid = '0' and rx_head /= rx_tail and b_pending = '0' then
                b_address <= rx_tail;
                b_en <= '1';
                b_pending <= '1';
            end if;
            if b_en = '0' then
                b_pending <= '0';
            end if;
             

            if (slot_req.io_address(8 downto 2) = slot_base) and (enabled = '1') then
                if slot_req.io_write='1' then
                    case slot_req.io_address(1 downto 0) is
                    when c_addr_data_register =>
                        tx_data <= slot_req.data;
                        tx_data_push <= '1';
                    when c_addr_status_register =>
                        soft_reset <= '1';
                    when c_addr_command_register =>
                        command <= slot_req.data;
                    when c_addr_control_register =>
                        control <= slot_req.data;
                    when others =>
                        null;
                    end case;
                elsif slot_req.io_read='1' then
                    case slot_req.io_address(1 downto 0) is
                    when c_addr_data_register =>
                        parity_err <= '0';
                        framing_err <= '0';
                        overrun_err <= '0';
                        rx_data_pull <= '1';
                    when c_addr_status_register =>
                        null;
                    when c_addr_command_register =>
                        null;
                    when c_addr_control_register =>
                        null;
                    when others =>
                        null;
                    end case;
                end if;
            end if;

            io_resp <= c_io_resp_init;
            if io_req.write='1' then
                io_resp.ack <= '1';
                case io_req.address(3 downto 0) is
                when c_reg_rx_head =>
                    rx_head <= unsigned(io_req.data);
                when c_reg_tx_tail =>
                    tx_tail <= unsigned(io_req.data);
                when others =>
                    null;
                end case;
            elsif io_req.read='1' then
                io_resp.ack <= '1';
                case io_req.address(3 downto 0) is
                when c_reg_rx_head =>
                    io_resp.data <= std_logic_vector(rx_head);
                when c_reg_rx_tail =>
                    io_resp.data <= std_logic_vector(rx_tail);
                when c_reg_tx_head =>
                    io_resp.data <= std_logic_vector(tx_head);
                when c_reg_tx_tail =>
                    io_resp.data <= std_logic_vector(tx_tail);
                when c_reg_control =>
                    io_resp.data <= control;
                when c_reg_command =>
                    io_resp.data <= command;
                when others =>
                    null;
                end case;
            end if;                     


            if tx_data_push_clr = '1' then
                tx_data_push <= '0';
                tx_head <= tx_head + 1;
            end if;
            if rx_data_push_clr = '1' then
                rx_data_push <= '0';
                rx_head <= rx_head + 1;
            end if;

            if reset = '1' then
                command <= X"02";
                control <= X"00";
                rx_head <= X"00";
                rx_tail <= X"00";
                tx_head <= X"00";
                tx_tail <= X"00";
            end if;
            if soft_reset = '1' then
                command(4 downto 0) <= "00010";
            end if;
        end if;
    end process;

    process(tx_data_push, tx_data, tx_head,
            rx_data_push, sys_rx_data, rx_head,
    begin
        en <= '0';
        we <= '0';
        wdata <= (others => 'X');
        address <= (others => 'X');
        
        tx_data_push_clr <= '0';
        
        if tx_data_push = '1' then
            address <= tx_head;
            wdata <= tx_data;
            en <= '1';
            we <= '1';
            tx_data_push_clr <= '1';    
        elsif rx_data_push = '1' then
            address <= rx_head;
            wdata <= sys_rx_data;
            en <= '1';
            we <= '1';
            rx_data_push_clr <= '1';    
        elsif rx_data_pull = '1' then
            

    -- first we split our I/O bus in max 4 ranges, of 2K each.
    i_split: entity work.io_bus_splitter
    generic map (
        g_range_lo  => 11,
        g_range_hi  => 12,
        g_ports     => 2 )
    port map (
        clock    => clock,
        
        req      => io_req,
        resp     => io_resp,
        
        reqs(0)  => io_req_regs,
        reqs(1)  => io_req_ram,
        
        resps(0) => io_resp_regs,
        resps(1) => io_resp_ram );


    process(clock)
    begin
        if rising_edge(clock) then
            io_ram_ack <= io_ram_en;
        end if;
    end process;
    io_ram_en        <= io_req_ram.read or io_req_ram.write;
    io_resp_ram.data <= X"00" when io_ram_ack='0' else io_ram_rdata;
    io_resp_ram.ack  <= io_ram_ack;
    
    i_ram: entity work.dpram
    generic map (
        g_width_bits            => 8,
        g_depth_bits            => 9,
        g_read_first_a          => false,
        g_read_first_b          => false,
        g_storage               => "block" )

    port map (
        a_clock                 => clock,
        a_address               => io_req_ram.address(10 downto 0),
        a_rdata                 => io_ram_rdata,
        a_wdata                 => io_req_ram.data,
        a_en                    => io_ram_en,
        a_we                    => io_req_ram.write,

        b_clock                 => clock,
        b_address               => b_address,
        b_rdata                 => b_rdata,
        b_wdata                 => b_wdata,
        b_en                    => b_en,
        b_we                    => b_we );

end architecture;
