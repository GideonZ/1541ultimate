��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]4*�U]'�an<�c�_=
N���G��/�G&,�*Ot.�+���ߐ8���94��s���r5�G;Qw�4����y�8����:و���G?=�XÉ��䫻G���c�����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�PJJ�6цZ?尢�e�k&Vo����?`��V����>H��=�e��U������ڏܼ�-����@������K.R4�t�Ƙq��G'��?�eg�� +P��W��-�׷Ypk�ݐC2%�[�v�0�-���U�_
g�>K�4��"g�XI�@|��铿����S%3������tc9�!�I�P�'���Mg����#z�]��V-0|U9�R]KS��Ą�>_�@����VwB{��=^�Ӂ���FĞ$[�k?�L-
�j��n*5�?�퀫����}y�W�K/����}:��A:n-h�<'Z����O���u�%����w�����bA�6�<�amc;�� ��'��a	U��-�S�d6+������/�e�<��I�ڍ�|�8�J���^�5�q{���fq���!z�`�%w4��沶YQ	�J����/��h�A��]���$����~�r�7�ࡎ�ߢ�����"3$s�G�?W����;�tX�%-���g�A�i�B�IU�p/W��3���yo<�[��\�le	�-/��Nx��$3G��Srg�A[���ӑA�̖���ǟ�L��VnM�@cp<,�K��:Ͽ�^v�\�1ݳ������g������ːy� N@Ä�h�Zۍ늩6#%��2 zH�Q��A�E�
ZjfC	�]���vB�����T���3��~}��l���@�K�Q�b䌘��@�ԗ���{ ����$2��J�y��5��}og+�>����>&h-��_�|�{R"-ؐ��Y|b�TH��tbz�U z�ƙ;@�@��LZ�M���Cxz�aq�W�y����j���w�L�y��C�U���������e���cau͏���"���O��r����'�BY�(:)d�V�,E$���i���]8�X��6�h��h���.DDz8���x�"D^ܙ�t}9��1��Ӝ�f�!���)/t�s*Y;=;��(��G�!�һ���(v&
Y���"�˥^�ډw��%�����A�m�B�rEo�>b�r��}��T�6�<�]�S�Ĭ�����S~'�����0�sCi�J�B�
�����r�]a�,���K}�y37���|���'-�,���.,���U��&�����/� Z�,�J�NI�U��ժ�����+��������/l�V�+�f#I[��4�>���z�yr�Pm�TXo"���@u�&��#��6��o92jҘ�M�* d���S��lDO�j��`:]^�8�����
��)g_E%t�$1��7D�瘁dW>�P��[ �fѫ3��z��֌ؔ�:�5h��ԲF�2te� ����^����!H�K�Jl��;ɟ�ֻ�#�s�l� ��]>:�%/Sj��.Z��]w�i�:قW+o���^��T\r��э��>���(N^�t��9�$x�
�H��|�DD'��-#�G����RK�]O���������[V�jr %�tMJ"��RWH2��g�7�!��<!��3�p��K{ҙ��1%M�������bu���u���Όɇ֞:�=�`�cr4y#4?�K�>�t�}h�!"N�X��=��@��[����ԊAN��Q���S	Rla8:F8�ngE�4_��k�oDÝ-�-g1�.&��y�B�W�)���S.��w�u�M.����I����p�*�6
[~��ڣG����	Y�q���%ПC�����Ԙ(��Ybפ�=�����JwY������!ka���]�yWm>^ȡ4��Psa�o2}-&���f:��Xނ�]�>9�'-���q�w�p�Ѳ��L���&� �}RI�7d�����i �B3ӆ�����V<1,I����J�,�	vTl�oxX�]����=, �!�ie�g?���v>q����1���N�%�c��/<���\!�dЯ������S�5�E*�V&�)g3-�z��zl��_��Bf�׶�Ɠܠ�Y`���!ӏ���L�g��S�`��R|]%$��M�n�3fov��%��i�ب�7	������J�����~���ʧ��\�4�q��}����*EtCVb��d�HB�o/!���^*[�� �Ť����������C���0Aҥ�}ȃ��tA�K D�=-C���u�xR����9Ԗ鞣���D39�O�K�|<Z)�?7�h �[�aX���e:<;~gD2C8^<��O�l�f�/1U�yp�wC@�h�,��YYD��*EU2�ƻ#�¶�:-�,����<Gp+��io��|���U�z����cn	�߱��IU�{��}��޳~b4�U�+yl��S�F��;*�щs�D;]�	��L+����]s.�<{?��P!@�1����ݱ|�W�,Uwu  �2���9�o8���"�Y��y�p�a2*/�Zl��lю`���	���ZT�1I�K�T�[I������O2��o�'%��b����\8`�)���!�^Z�懿�T~܅g<M�luˁ�R�LQd��"�$_�3� ~Z�)Hc2k�&C8�E@�鵞�>��P���l~ܶ��v���� b���(k�V��i�c�b�ELV�q�`҈P̙y��#LS�:�#L�U�U��*�?�R�q�N�+:|HMV�C�0-E��1�[N�ޫ���WS����B&@m3�-���{�Ä=k�`ڲSx�˧�k�W������_ ��Ƕ�mh���@�J!0�� ٪�Ȥ7'����Mw��|�vD?�w�QCe���[ԖЄ`�G���W��q��Q���YgX�H�#���Ƴ>ɵ�kH�H����˃<�r6݄��A6({:��Q�o-��urD��'������f0�ā�_�	�����E���!�����{$��z����U
 �ǵ�گ�����W�phhmEl���I[������e��C�<h q¹���_����8_4"t��u/=dxvpQ���HM���&<�����%��G �C�Eb|p�.u���w0��-oW���lj�������9�E��i5p�d�1����:I�B�,�D��t��>ʭx�E��5��-��ڈ���<K���	�ou���1~��Ӥ�T}���vw�*^ ���=f��O(m��n�D#EV��Z���Vxa9hfj؀�D(��0nO<|���h��(���TP�6&�>@��	�L��WP0����ᵾ��� �{�a���
��M�бǊ�&��?$[�4J '��@Zm�(��4V�"�-f�7���U:k��N<kw+G��/!
/���'B����T�;�mwC�|
m��*h~٫��|��q}7?������Pc��)��ѩ��g�4zt���4��'��5���+CR%�JC.�C�_�?Қ�;�����#æ������v)Y��^��fo?vMY0��,V��zCU�A����e�ݦ͓7C:���
�>�2����eX�X���$��ZM$t}t�!�v|��ϣ��N�
ӹV
�\���^��R� ;��&�;���NМj!Z��חf3t�H䕭����0�B��l��a9��v|�����[GyI��������������c�v�^����*qBa	j#M��zԣ�z��g�w+���IFԑ2��wC�������S��*𐩮����@v�ߎ���V�_��J~������2�NeG�W@����'�'�Ao���ϰHȥ_�RJ�`V��:�* N`��a4I#!����g��T��4�B��x ���rceѐ�2��@�.�$*���rI�ml���=}���y�-���kЊ[P�
]7_��h/�O�N����/JyNx���iE�ފ���>��NH�
)gS�r�y�0�G����8X�%-�"��M]`�l�0��[Ⱥ�.�~��>5�	�]^�J��G��-^��[������苖ʎ�剷�b����;w���|�Ʃ0��=�ڐ�0��TϽ�ѝ�k���+�H�c�0ʨ����rn3��a��f�lE��}\�mQN�9^�?G8v	��q�4�O�*U~\��h� ����'�F��M�9�*NE���b^��9���z	���k�����X4��r*�xVk3��Qd����d��Ɩ-/$`����R�6]	d א�M����c��{z�^��Y����5�\:ؠ�Ѩf��ji�� �(��t+"�2ӄ����1��8��ӹ�r��ߐ�b�e����yE����g �ȍ0�:V�
��*�at�� ��q��q���p�lv���z�f�T�:N~�L���h��:�m��7���*���a�*�|�V<���\$z
l�8xf+ȵ��e�0�7�ȱ�u�̎̏�*tx<}�&��Vv:��N��c~M��H�8h�,@��G�:�Z�[����Dƈ�d?Pb�p""�.U'N_��)�3b/�P~ƞo�@(���� �C _��;������qN��PV)D�Wi�}Qg�2��C,��Hw����@��RJ� L�
��=0*�q����x��Ex���K������]�X��m�y�|^6}��P-�_����>�Cv��'���:�%���"3�GUN���d!
�I�0����pi��t�g"7p�c��f@4<yyR�0EK�怶(��P�@�t葸L�!��*gb��	�2J���. 2l�Qv� 5�~FؤeÙ�.㢹A9�(!]'��R>+����*;���4����ɢ����ȭ�8D'�!w�X"�K߻G�}�:Ɏ���ɐ����]k��-[B�z�{���4G�SA�OE�®yF�(�H�hI��zD'�7��Zx,������3�;���H��[�	�.�6�ՏkKџ�/�&��ٟ�Na<��6�F-b�0&#���]����g}����\����5��������eQ[р��=��s�b�Vx���Gp��a��q���l��;!����M��!������"����$�F��� s�P9a�܎�}֑�UVRy���Xsj�x��Wh�����!�-:|����h9?�|�/���$㼕9�����^no]`ʷ�I��%���N�(�9�`�󞧣,a��.�-�:����v�H�?�O�"��L����H= �>d�&��O�/��kS
{��q��Ԏ�AT�s�^�m�;��7(�.-[��mnk�!�>���p����?����R�d�FX臈[>���M�֨�}!�-����#CQ�mn� �H5�b��y�Yop0�a=9NA;X��c[���;BՊ�h�1�۬T�y͟�#}�1�6#G.����DV,��N�@�XD����� �r��{곌ih�tT�4�e �i�A�I��e
�>$6���2a߈��K��y����pQ�{�Vc��3ѻ< ��D�q��Յ)�c�LB'�4f~_�_�%�3rD��ᷧt�y���p�ae.Tv ����P���Gk��v@P-D�U*��
�����{=3h4������s�1�c��|4�U,�9ȵC�.ƥp��4�s�t��b~m� �Ar����l���H8�����MV5X+0U�̸�C�|��RY.f8���� Z�>v]���b=�o�̩���xCey6�Ï�1���
��b���A�p��������}�|����#�͹��[�š���w7�v�d���/�����B�b
�d���n�N:�X��rG�8�K"���\�xv�I�������"�P�o��r��.YF9���C5ץ���h�GD��������>$�	�|�,����t�8�o]������,0�$ש:"W�<���L"�v�8 H�4�F�~Z�E=��a�bCJ�w�{�s �\��M]��e�����*Ӽ]2���R�i�J�u���l��؛pS�is-�;�0�p�na,���^��r��uG�?q�ѻ9b@��7��c�xiU���C�v�ÛE��&=��&��Lx���rA>0��l"�p�#Ѽ"/r�la_��b����F3�TsP��K�m���$����P�<GX���9#k��xgܹ~���9t�������]��k�,d����j���-S>?6�,G,���&⣌�`�b*_�ɼ��|�­X�h�b��NgX�o9=S@��Ǟ��x/P62���|D��q30�ו��9C�fm۔gF�Ģt~�}��b`O��X�>���A��sO�/�K+8���G��Bͅ��Ԟ�%���fs��9��i�����z+Y�谞`�=�I���y	���H�whHgY�M+�T�����O-OesR���t��j�5<ɵ#/�;�V �_�*0ua/���	�����Fw�����f�U<�Ε?<Mxk�0�s��4I��]~��%=M���&��Ǹ��O�٬���p �����D'Y�ݪ?��|�=B<(r�X��nLϽ:��(�$���$*��eFG~?�<d�4kz����h�-��Q�Q����&�$�k�\bT.�.<�η���u	g�r����ʭb�|�Z�"��f����D�,�
]g*�ZN��̈|���ځ,��'Q�!W)m��ܗ i	VO��5:�� ����&8�^�Ĩ� ��&��I��.@G�! RŇ�3�Ӝ�5=_��˶~g�c[�F��l��zӧ�r��=]"���ș�N:�:S���L�';e���	0S�����2��� W/giG�q�I򕞇 ���d�Q�[���o���Ɏ�����)����/������G��SՅBB��[`���>~����(ܤ�m��VKl����" 瑌xD�{\����`Q�c��OϤ�Ì����o�	�=����,[�f�2)R��	?�c=��63,��"�~����&):��M�譌*�DF*8Z��ϦQ�=�Yj�!�o��MIN�����^���o4�:%U�=ݠE�{���j�:,�Aό2OHA�"+��)Z��`χj���4P���^�|GĆ�M̢����I�y���*�GwR����̆;5�ڂs��+��[A�T�v
q@1*��R�+Oլg�t�����9]���c��%�`�x���ֻE��g�V,�`�鼭f���+͎�M^t��X
)ϔ\+�z�Y����:Ӿ��A�Iaͱ �L>��������N	]���~<i���(SMgIL�_1�J��X�|Ȭ����9K�m�\-V9�*����$�fq�������da�E7�bw��~~�(���^���b���.���+smBv-W��P����a��:)}���**^zA�6��C)�I8J(��%�������['�Wq�B�/H�Ywn�4��{��-�r9mL��O- E$���GƑ���X��E�QX�|�#]��6���!Xk��$�?(K(�����Ȋ�y�6��\�oy0�d�GHS1�y+j��8��["w
�$
?4kˇzw�V+j��}�U��� v̽��u�.`����u��X�<$��̳��b�������f0�p�c�u�Q�F~�j��5�X_��h��]����ba������`�81�&���_=̗78��F	~�'S�h�+��K�;�q�u�b�7?�-'0P�̍?/��۴RE"ҫ	�u�"�}U/��r4x�N�1�_<5�%b��B���f��A��D��ד��v�SYW�/eC9|�*����3K;U	k��@Z1�"s�}D[~�Ye� Y��s����-��LT�ty�dspY߉ 1o�ԃl��2p�/'zBt7yia�,S�v��c5ݿT�'
�,��.�o�2Ⱋ64�
Ko��d�������!R�l�b��7婷|nU�����2E#/��0TY��0p�˴���1��E����������I�~�<cv�4���Z�A��d�fY{��C �e��o	�N���(�M�uL!�K���T�f9�|����1��mA5����E��m��8�B����6vmF3�I�'��p.Z�։�Y�36z��/h�.Q�$��`�p�̚x�����Š�QXTa3V�����k� j8^t�u����8BW���z�r�%��p���g
SU�,^�Ԃ����#�"�ai�^e�f=�r�CF����>Ze9���|&?�_��J��V3#�ٹ=��&�:�1��J�A�_A�I�G������ѹu��������+�4q)��lୁ�+�)o��?�� ���u�J\��*x{y2�P��%�f���6�+����2��'���_��t��<��&�%n<�*9�;�[.NV�w*CC�Ukrx�gݴK3#9܄�ld�_��q�.�w�e�,��E��mv�`,�R���T���0�ۥ ���&�]7��ߏ��Q��j�A�Vc?�#�x�� �C��?3�<>4�S�f��,�Bi#@`O�3�:�,B5N�F�I���h������n)���\�W��;�.<�%������࠙5�����KΝ�����vJ���5�+�	��&;���)���ʺ�&�9�a���J�c�����Y�a��r�hq��xt�
My@+���?���ft�T��6�{{�h�p*H��q���3�U�(�!T��(C�pG�ء?7�b���}'s�!$�v>]�����d�|2�6��+Wլܫ낃��R�"Y��D�=�T���f>Z1��+7�l�n�d�����M�#�����42z�x��s�R��y`%*ߣ>X1��!oO����������-����;u���-T��QΛ����%���ë��b#a��r�ػza����'ݗ8��Z>5n�w*n^��׊�- �oF1Q��_j ��0M��;	枴6~0X���W�.Qŭ�=��<��lMM��s�\�ޙ�o�~�	�Q3�48��2`�+���X�K��-��GW"�Q�D|m�n_�W��L9?���ǒbc�B��D��q�`������p���-�F@[uu{{M�VAJ��N�߱������_�/r#��n4�g#1�B�dL6ۉ5�|�W���/�'z�M� �aW���%��hXԊ�����TkSP��������'yG��zZ
�жh�]�s�6�8�m}�#����7���q)VG�!�2[ԉ���	���#���.��¹�m�����R�C|�܃�c^,�V�9�LW�f�����>8�y���Эm8!��2Ax��_v�Е-Jd�\
�x)��)>����R��|�w!1�R�J�*���hM��"�,)FF*�ۡ�J�M�p��Y$�)"�|��,&��ڤ͐�i�4v�Ņ��`���b9՝�nVxg�S6����)�L�A^e\�q��ل�7]������S��my�{$�rG�GI��&} �����
n�\U�T-��G�=T�DY�k�-j������6�r���<�]����fJ�p_ h|7�	�/),�^~�	�R�
�K� $��q-,�c06��,�m8^��7;�]��~�����A��qu�ǅs*��u[���yPpN�ӽ2��>�5(Jc܄��x�!�9
��mq�E9"\?�>��!>�����8�X� ���y�k^��Q��C�{�)D�pnc9aO�V��k"��X:�}}V�_p�Xj;;z(��(�.��n�$@e��zm~ou_�l�0��4_(�{����w� ��,/.*�Qe�\�LDɅ�=�Ӏ���3b��5�h60�
��?۩Z�/^6��$e9"�5��`�D�Od�I�('��L�gdfS0v�Ħ���Eb��*>��PK��I�6.�ƵS�đ)ݒ�t�tӨɼz�Q����Z?7�̣�������OE��]pDR$���k����?Ͷ�K�#;�9�k��"��=�.'�P*՚j�x�K�؋s�Mk���Ӭ�!_��StBa)�E�ǿUp������\�y�]ʑ«oN[֯�I�t�u�+d��el�f]�o!��[��4���6��n�k7Y�o�P����,*]A��D��B��g��cS U璱#	t8$�&~�߰�����G�{8_�>ke�����:�H�.��*(���ۤ�� ���B5oe�Q�����t�z���栗��<�3� J���Zd=��n�k�@fr:+}qj��uk ���G��0�S�����vLm��z��8j�{��dyI�9�c,�^�6���r-�K��lh�[��e��~�ޞ��Fp�,�?��l��@���}AH���f��5����b�º�Ȫ�T�"��9�n��-E�Nx&���k��&P��U��oVa���Xi���C�$�+BM�Al�my������L�D�t�D�CDF� ̎-ot�����",7�Y�no����Ca�
�n����Eؕ7^mb�9@����@%p�v��oYf2-��Pl��ֻ)ӹ��mO&a�5,IY=��٠���Ha��ٱP/H�����>�L9���R��:��������ڢl�)D�v��C��";W(تd�]V�~�t�H�mc�B(8	D���~S�ŏ��P��ՄL����CR�$���<-��k�n���<_�v��͂2і��{[vi7��+�0,���� ��$�C�X�9-��|&�eٛ�Hoz��;�[���Mp�	h���\k�9��P�mƝX�I�T;qu�>+˄$9Q,ʿ{,�L�n��I�V+M�g(w�]���a��*v�	Д���ۿ�i��L�n~���I3y��'��ޖ�e�u�#��+�c�IS*vq��j�Si�`p�W^	dK<�!���ۊ�d�o��e���$tM�W:M��Ym/��"Y���y�i��J�Y�E���Y�b��_��7����a~�s���{�LK�����#�F��,����lf�6٘'0-d*Q���/D���Ȗ*��ȠG3�/:����e�b0��ow�j�b�;� 1r���Jq�hE7��RV����m�������$��w+���mY������ CG��Yܞӭ���)Ph�vmO �l�4��cEK:��!cx;s�<����~�|4�Y�{�p�<����[E(h�Θe-�Q���l�4_�״�2T@�ʝ������׾���೦'%���X]J`�����O;�ؚ�8��r,�k!7o:��E�Ӝ�}I�5~� F�Vrg��ٜ��̔���Q��W*�3���3���R��ޝQO69X�\6��T��SBR��,p8���S�=;el!q�h �n�[�K�धj��e�hWRƎ��"1f�M)�OC�F�f����,ۓ��H�3�;>�?�U3�0_.�������S�xc�Q坐?�X7 w�⮘a�ʿyy�%�W��z�E�Kr��]�ls��0� A31c�A|��w���������u�v_���l.@�c��2�>��a�eH�_B��F�VK�w�Up�@���2�c�<R��Y����l/�W��q\��#�>�"Wi�9�G>�=�aD�����87$��w��%����[��>y6%�,�t�D�b��ݹ�5�|��L1s��Oe�e]$��zP0���a�O��_Fܶ�5|Ӄ��$�ݘ�L��W�@0(`��������,]�����r�й�?��6��C��x2��۵�e��:%rNxN!𝾨��Il���s���{N �t��ջ+1D�r���@YN�ڿ��6	`�&2F^���) ���yc�z[��ٗ�u��u�󕏕mB�@���<�G+`�9�ψ���]�
)T1�����=6����{�T�@�=���nOk��퐌��vK��}f��xa�h��k����B�~nNJI�/"�����b_�4D�q����Q��!1]�v�,<ӯ�mة�=�G���7s�f�܆���5���1p�W8Lģƛx��^n���=�G��^viErW���w�o�٤� �J/�ݖ�y�չ����Z�xYx����Ɓ�
��a�{�y��`���-�(a<̀�NzK�@�E �����6�?/9�]T������o��N"��X�N���b��S�SL�J� <F.%^�X?�J�9j��u�����@&���������E���2?i��o���Q�9�y�l�X���bA�\�ћ�C �As��9z���r�c��F��^Vф�q!�r´�xV�́Z�U^�C�Y��*o�.��< Z؝���'�,�dz��]Ru�)��D0VR�x��s�J�-=k�,�x�$Q��+����WG��t�);�������V�N���_F�Q}�=A��[#�h�tg�ޮ��<2�h��n���q��mk�d�$��O�B�%�5P'h1�i\�^:��Ld��9���b��X�H<p��<�Ƴ�{����w��G׊|6���O�ܻ��v�Nyu����c��#����]jA����y��VI���=Pa�x�z���b�oX]�ecD���4��ym��D#�*C�q��J����9)� �ax�@/7/�,"NsFy,^�PY\���ϋQIĸnڟ//,6��(]�m�h����R�K,�l�W��K�>h�v{�0��d~�_Vm��D����G�e�'�������pß�a�ݙ����A��-6�ʅ�:�
���fJ[`��|{������=�y�)=CiOf%�e���6���kX��^:G���k[1�-�%��V���"DQ2;��)����:�%?f��A��}�؜�ƈ[�E�BZ�dl��t���6f*F�+X�J���{"�����|�)��G��H�`٘3��"V6?l�L�fZ��@� Dٲ[��5����kk���,į��\�d�)u-��|�L�@0t�c��x4�J��V��%�uD)�œ��$i�U�������L��#w1[�{d����:��'AG_�;��c �8;�	��6m��87�8��%����A&��:\,�F?��`G�1�|i�>�'ǆ5���MƑ'�m��7�^�6���w����kDϛ�}rvb��avg��xnr^���KUQX�a�M>(�*��hFp64V��ܠsk���LmW@���H�����J���b���:p�˧�IZ�oH_�k��ײ:�wu����{{���a[-IP���q�a���.�����}���ϊ"�B��;ء�x�pYH�짉E�b�2�Ӛ�0H��@8���.Y�!������}&f��Yb�����٤�߼H��A,��&�1�䂴�Ȕ�Í�͜��>\6��jEn��r$�%���~X������J��J���$d/XZ̀$�O^#û��k��|�0����nO��^0�t�dҪԯ��B��Y�FGJу2!�̛h{ҳ��A���.�Mt�yϋ�Sq�����eB�XcCZ�`8*o�Tz�íX����Ag����b�E���$T���o�G	��^R��Vެ~AȠ���瑮:~7�&������R?0|/��P�VL�S}�s������`�h3�R b;��O�t�:�?�ð��(-���l���뷹���V&�m
:��(s��6�ǔ��"p)��rL}��[�!��L.{�/��*�������I��hx��B���!�+ Z�S����{ܳ��e󩅝��{�^��;L$$gb�6j� ��2�.n�X��@$�j@o��;�+kH��ۦ�)�
�3q�Ղ5אx5�iy�'c��>>�r��FV���~q*%�q�ܧ{����䂓��H$�XZ���?(�1��	q���ޖQ.w����Y�[�	2*�� L7d>���w`S�C�2�����F�Y^^-"rv�����K�3�rb��!��	C1I�G�f�n5��`�|�8�bC�ugoD�-��4|k^*�	nΆ[
�7eo��H2E�yu6"�t�G�`���`�t�Zm"�]+��[����8����F(Mi���r���)k��)1�$�{lowcnx.�Z\�Z��F�Wx|, ��#Wn�̬��K6�6�`E+bѧ�$�>�g36�/��|�<�\5�rk����@����4y*p[-��4��c�|*^@��
!�ʒ��Oz@74�R<��q�Uʨ\�k�U�T�O��8�5f�^��������՚H�e�G���۾ΰ8Usg(�	R��M��ad��v�\��gU��|�*y�C�z��"�5"I8K4�zE�"��Fd�4��"����#��"榾~O3i�����ABK�q�k��)�*������/9{�u�hN-����M���ą8��i��9��c��ڍ\�ް{��NP|�E�I�����뙀ݐ�	�����>P7�*��3�>�nިa� �����M��u���;=���LZ�+<M�,/N�y�_R4z��!t�mnw�ȑ,�Z�����2���?��m�j�yh0�v�Ļ�<���=Qne_��dքbg�h��l,�|�����o�Ƚ��uf�D��Q-�E@
� ۧ�4�^[/���K3�U�p��&l?,@���8�e��[��!&��k[XW�t��w�x!�=���)'Xj���ƕ�����>�����//�i�0Ch�#P`�����FT�D�PG�|2y���.b���7Z�&��������7�}�kY��0V�*����J��?)�'k� ��v��u#�Ex�3V+~�¸ �8ۚ����	�=�	?^�o��/JVIm*l=x_%G9�o��i�mY*�UJ?=����h�^|"��=���WR�!��1f!)������7�O��hĐSZX�-P��"e��xOr�d��K*����!e��X����g?(_6ǻ�!�T���W��oQͭk��ǯ"�"�����3v�K+��~>!#�=dOܚ����K����/�M��.��5����q!N�u�hO��O�(�X,7�W$RKF����h
��߰��P~�'���R�a����TeQ��J��h�<%l�E���ڨ�+��fA~�o�n#oyw�r�0]+����q���S|�ե��RD��`s�������j}2lZ`1@ms��B䢹�mҢ��S��7��x��軩q���Y/Y[�w�B�4a����F���j�]~C8�uG��F�� ��<Pו���1��.�X�� 0�j-h�^���RߦB:�/��*��*U���-����.eea�Ć�w<[�S�W�v/	�q��L�y�w*;��_둠yӫQw��E�-���*���/��;6M������x���#�Cuָ�A�$��SeB�̦�U�m�\���^J����y�J��l���!�v��o_�f`�ȤY�Ȳ �"��Rx7S]څ�w�JE���y���)��x��w�B��s��iq��*����P���	��B���p�}���Oq�+��	�ѥ�p[��L�L<�N.;�]/Y!�ҩ�k|�E�e@.[+�FE_�:x%���{�Nh�_H辿_�O�w5�{�$����Ү�������T�IJ$��x<���ΥJ�\�c�zm)�	paK�>��}6V<��βܒV�s @2�:K��r��f(�38���S�\X�

��J��3pC�-#tV�4Os=$o#W!�����Ov�,jqĐ���5�G������)��`�G1��J�j�'�����x���]NV�L���C1Z���i��%EXSxD�j&��� eɚ�'P ���h[���wjW�8��� U:�+E0��t�Y���MѶ��"��0
��m�ݲ�� �&�/aq�1��`�F%p��ͻXd�"&A�	����
iΦ�C�][�A�vn�kˑ2&]����Qŕ,�&MS��n��h���4}�[d��W9�����k��$MH��Z��!�۪̿W��_�����f��h��QQ����s���<�f�����������в����I�(QA�*S2'��#���H��F'�Cr_{VY<Sp������0�=:� o�|Y�	c���)��	E)O���?�Fa{�r]�1(�R+�1��(W4�)o������~$��Ux�S-&b��!LP���f�ݗ�<�p�W5�'|&������7��hd������7�IqQ!��e� �#YH�r9�p�%�.LE߀��f�A�>;��r�jD�U�1N٫����a'�=91�8�Ƞ�A��\Ӳ�=���$�bT��� �ىY�1Z�,�`�cѠC�u�I�Y`�Ѝ� �Mp��/�K��\�I�~��|qS��`[X)�Ý��O�4�ϦJ=���/�d�f���
���{gl�ED�H,����D�N��@�oz��_QDn(V��?O
Q����*1c�)4ީ����:h��6@�RJ�H`�%"�"/@�ט���RD�n���S'�Wnj�����f�gU�d�ObX���D.�}ݲ/�2Xo{��?q�j����;Fx! �	�����5��� �B��D�\llk���]����2�_�e~-�&Go����Pty�F��\��g�w-W�(���q��7D~��	5�(��^Ý��=a��m�?�ύ�ꍞ<�8 �m�硷{NBF���>�+9b'�jnN̩��+lȥ��u���ǆ���U	�#��*Q��w��{񇾾x3U�	�̽�Q"#�F�hݑDy +g�5z�Zr�-p� !��p>��C��:�VT"$�[�"6�c>��C@�+\���XL��6��B
��3����PV�4��&Ӭ斛�^CM�Y+���Us�kQ��лg-[?�t�Ɨ�<�����R���I/�}d���#B5��$��D@�l��	N^єHD���D�Td�ϝ�q�^�3�������<'C&��|*J�3���������ҞK��&�ǌ��o��v����;�	-�6�:�v7{B��4~�8w�N��BoF��>Y3��_6��E�!gF�+",]�]Pq�%���E�;_�dZj�|��b���AO% ����χצ��?zx3l;�� ���,�}������.�w2Bu|co[�b
�h��fo��<Es#s���D��u>)��U��Y9Ϻ��+�Z��;j��	7�� Q}c�v\/�C:<1�УEx�Pp��ZN��Z��[�z	svڧ�'so��p^-(���qjc�Jfr|z�iǻ6�M��$��/��,�@��y�.����Ѿ�Ӄ��N�,d-/$�:&�A�-�8�zT��ȈB�k;=b���&D��k�����)�p��+�Ti��6�raW��?�(ݸ�{��6�%9,��G���<h�:^��h+O��7�)#~�>�����WٿMܴ�l%a�Q��$o8�s�`�Øbv�jm_�����h�:�<�����MO�|���βI��{l��{v�T�NY��;�T�������鏝�7eԲ�-�д���!�܃)��=�q�d��%����&���,]��r�uWV*�4'D��8��S���kأ�qC�|<��:K*]�J���[d��'=�)�z�8RƔ�n�-:��!1���f0��z��(�6��O0��2*{�ث��ĉ���O!��]�a���:D�&���LTL���O��Y�	��6~�D��'���j�
��Hϛ3�_oF޿�-JL �X2����W���"ˍ�'\�
����$(��������l������MNd����k�h��)%�e��=���ٸ��$�N`,�'��1���Bg��!8p��,&�s*7�p~�<*X@����$�w~��B���x��]q���TV�^��*�;X�T��P��gJ��b�����Ǚ���mۗ~0���yʩr�.�"^��NO�����^�#T@��74/1��[�d��aH��\E=אָ.��u���gm��Q7�Qi7&pH�I�:z�k��ճ7�r�/F�!!ĝ ��.Av
9�糠��췵��*~Gޒ�?��'sz��a,��m"�����g#d��{�萬g#!�����Dʱ�5&%H̃iƓj=�]G��"��;��L[�b:s�,�ْx	"{�Z%.�>���ݖB�5�kdP#<O��YA����$4rE�VȮQT�j��VtԓMZ�.���&�&�PِM�}�ːt���Ib?�R��	�	�V���4�H�L'���2��Q+��g�rN�O��//��<.�u�xdA�b��1���+��L�	)��^�x�����y~� ���a���q�i�AZUVE݅������]���B~�;�K����(�e�Q>L�c_{5�F;�b\�d9��p3�g���[��s�G��]��Uw3��U\n ���C݂�tCJ'
�ea/Fk�T�̂���c.���J�bN�w�8'�GVt&��x�Y1=J��~,�`�t��=����Σ�B9���N]��,e�X��=mFFjTe�ߚ�]αJ*cL�O�;]"6R v��~,�F���\j*�#@���t��X�$�;	�(P�=^j��y�D���>B�,��U���W�!���
q���cj�H��Ygʓо��ē-¾ٚV~�?oL�8�4����t�?�����ܖtŨ9�a�-�e\�����������Rɓw���:P�:e�!�H�>��ĕ�i��ֿ;���T����O ݟ�*'.�^tSzl�sp+Y�_�ƶ��W�i5KK7�!����!g'4���Vi�}p��Fy��{9n)��8��K���� �et�@�I��Z5%�t��mi�o�G�Y�ܡ2�X��Ep�F��GIf"XJ������ w"���/Ct!"�`�wNj;������=vE�I�ؚa��&�k[����]MsO��}���loviF�G�zV���/�����&O�fC�tBat�캴���vy��#D���[�����Xr�u��&�����`��1�&[��ir�Lr3;�^-qRk/4�\����M�JU���+uv����|`��������з6�?bǶ0e;C߰�&�1�.6�������#�p ���w�E��e�KKXۄHO
�|6�ڏCngG|���<M�0�����;����M D!^���S�U�a��p���,��vֽv#e$2�P�pn�u�����<�� �`G9����u
b��Ռ���`2�-}r�,D��#����XG q�H��ٿ��z��wle�4Z_( ���Y�䶁퉍��BN3Ș�f�>�幪�N �����B��,&��r��X��,Kr����^�|�#ǄY��l�΋ط�����tlQob�K���n��Z�bnh�e]�	�}4]�y�p0��	�����'qc�j�*�gU�`"�G�
�{�_�k�+��N�o��S����j�m�����
�T�gܘUlna���=�g���73�L|����NFB�۹�[d��P��V� �\�a��W'�%�	���H?�+�-f�!%�^���UUI5,nf�¸�j���+`��5�tA��v@���ٵ�~`8��+��Kl=e%
���]ǓQ������nwq˓��z�dv��u_�8�o�S4�@)_�4T{B/��2�%2���w����y�zX?�ϾpW[*߂Oi9���N���y���vA��#�+x�t����G$�g#,�����7���_^�$���p���J�u<����`	���N�P|�(�i�$�M2�B�����ͱU�]`ܹ*��HsI�����nI�1P}�/���)����
x����8ą$�1�9K�������4���BGNGٔ]�!:.V�r[�p�?�/Gπ�{3꣇�@��ѯ0�
����w!��4�e�e6D��k�������>P��:�O9�,���Y�s�xl�+��.��9 k�x2�t+�%}]�lQL�\s�0.�5��W��:�[l�z��`J�6m����C�Q��pY�$Q�K�I�9�?�� /�4+d;l����rxM(�J۱Zp`pI$r�޲xc���]I,�)���n~a-f���k�4�w��-�D�]7�g�~#.7�#v���ه��qt�0�Jw]�<K��m1��A��t�Q�������?$nhoR��'D��^����G��eO�"�S���2�����(!r���zyv�?��m�	��8�8��&>�iQؒG�+Vzv_��汒Wjf�%Ҍ��B�d���N.�b*�JB��N��T�����r�i����B�r��l��Z�k�j�N�l�h5�5{j	�Cl�}�_��>�pZɚ~�Tj���o�W���cr����FA�
i�Jz�@����$��X�^����f�45���߸B���^@Eڲ�he<h&Y�"�{�-�,3�_#4�t��'EE=}�()��h}h������e��z�*��A� �������I�jTu[(�l�~�3�sn�U���@cDfƸ�����x�).J3�{��;�33�r��כ���o���ԛ�z�ك��6u�#�r���Mm��Tߦø��m�+����E'q�,$���g�Ɣ�X����"m����zB��W��?���Ӧj�rdx�������c�+��L>���BV�+A2/f2�6"��_:�vK�9��[�6h~ϊ�ę��me��_��Pj&:�?��_;�͢蠘�y\�mn!3fͼô>�?�uY����m�m�DM[���9y~��h��)}V1B%�>��4Z��ЇT έ��$��z�Y�y���9�a�<����N:u�<�m0����� ��!K�0,���D��yOR��^����tۤD��u����M�,N_?�D[�
[-�.�X*�$�[��5���6�@3G]wɦ^S�څ�{�Z�z@6wD?��qV�/���I�7dx�;��d�P��ڿ�Vܒر�?��uJ"�
�st�d��&�Yv���V۰ࢼ�*��Dm�}��D���F���~ 3����Ӯ�qUi~YƸ�+�4���7�g�j�a������b�g�Pf��q˨��lr5����^�Z�K|��az~����l꘶>>���~�I�ӎ��4��k{?h¼�¹���?�rr&��P5�n�� c���!�f�M�j�=�:ڀ5��w��faX�=��ūmDgf	�G<L�f���acvN�)�o>��1��>�,��.p��y��?�i�9\duU0z�HH�m0M'�fE�Xlp_n����ˣ����|$�\��T(�<��������7{#+��<����o�z_�����s�������%�w�AlΎ��T�i�e=�j{����54�b�Q&��;�w�u�O�~IfS'0��~���Bg�Ԡ}��ӦݜZr$�U���tn�����˗dً�!ذ�^�9ʃfQ�p�o����䥆|F{�$��X�K���Os�^�1���c�y�mP�7긒��GFیޔ�֜(FEӘA�����q~uX�9A��.!���	k�=N��]!�Y{�S��S�t|�xn�ݳe���Ou�eO8/g3x��$�+�B��!vDd��7����M7��� x<��b��t���X�/����G@+�y	�;�z^���u)M���kن�FV2j=?xJUL��P�C�֒����݆������͞�W2Ո﮲bʴ:R��Ԭ~ �F���LN&E�i���*k�dֶ);��.ac�(���R�\,��cc*����Z���G��oJ����G>���51}�'�,|b|[&��^�9LA�d� �+���f��ٖ���D��R"�T+�C����� ��Ѫ�$Rf��k����3�1iy��%�Ø�#�d#�c����D%\���%���>t�E��?W�O�c�)��#��-��8����\�)���H�!��B������%�f��{����p��9��P mb�1�g�����ȹ��"=���-� t��/�Ia��t���c0
�X%�|2�ۈ�O�)4�tC�nA�h�aɏeh�2��'�>=@�t�}A�{����^5/)H.֍��}_h3���� �t+$�z���Rs�g�L�栃]���{���j&"E'���?�r�z��6=,Do
ay����4� S�K]I rE�d�Ԍ,���aG<\M�f�Ǝa�)�1��'��cPo��!o(@O5:���`Y8�|˖��j��������-2b�E"�]�Ue�7������ARo��T��h9��)���~R�Y��-x�@�c����O���c#����"Bv`�[�V�-n	��kH=�TP��fᚈ�}T��D5ɸ��X�k���l �G��4׊L<H�j�B� d:p�i���:Wf.�����w~�p��&ZȲ\#Eͪ�!�ź�-r��
,eЁK���)��-��u�	.R��J&X�� (��6B3B4�Z��Ҝm����	����-�x��q�V�ﮬD���V:zF������Î�;�8FIՉЃ��@��j�	��#���LB�E�:Q�aw��^g_�*uP��f5ܘ{76nHL���1�	<��������jv��D�c&�hd��1����*�����4sMt�H��?13�ߴKH�0Zq��*9g=��͕��c\7!i��?�z-�8�*?�yE�FY��k����x��x������'$hur�M@���\T�M��V4��^���!�x2�Ю��^�Rep%�2��k�uE�� �-�y�Z�+pӋT���0���~:x�0����nr֙�(̫���.�b����>�&��7�<BU�7�I��m���{���9��S�����$���Yt6����׊
	���`�s��p��ꃙ>������7.�N��%�T$��?)+�m��~�Ϋ�d�YJS,9����/�{/W�Y!]:]�'7*�4�=nI��Na����M�2@F,z��$�֪1ʑ/�.�F���UK�8��&�81�s�{���ƤE��S���>���p�2�q�C���y�R�[d�����`����B�[�{},,���!�!�t��&���&� ��[u����*��5�nBi�ŉ�5q���ɘ��q�|�|�<u������p���� k6�����|48ɪ��n�-�]������φRa��k"ˎ�v���>�X[Z�U}H(������ ��*1��Z�-z��oT\��U�>��EL�Bu�c��F؝��\�ع��& ����}z��K��ʲ��=��mX���wb����5���/(*�]@��qҕ�F$'S�O�+�Ӡ�o��N�^�Zҥ��A���6�T;T�"�t�T��=\Ήr&m�,!9c�1��������9����뻉�lC��:z�I�݅�;���T�S�	��i]hL岱�)S���/��!����f��#�E�tF���[�+��E�-�uD�ZG7�V��Б&���_x(���?_�V'�&�Xk�qf�u�����e6ϙ��9w]��!��q����@*P��G�ʶ�AJ�69��$�)j���׫�N��Z0��՚ϊ'5�D���X�Xe��.���G
�"3pdJU<D�/��'f�e�0$�WFjt����r%��a �c�� �ve��n����"�1e۬�y|�t�U�Q�xт��-���8�>��:`����;Jj�q��[/�K�tOUWn]�o>[�n���.�l"�U(.H�]h5� ��??�A[a�������tx�ޤ$�kDC��8:?�� �szPHe�Ǻ9�?��*Wn=><�K�QL�����������S�ˋY8��_}��E�/G���������Mm�0�s=�� ��5G)�X�>�������C��
�z�߄�T蔷ұ��]��PM��6�R�-"ײ��3������i��Z�S3hs�Qe����<��� "9�p��@I/��7b-��l��]3,�ٗV����	w3� ��;���V�p��U�,֣lD�Z=�g�+�
.�2����:���mC|�h �j�@�0�hW����Ϻs��0!yDJ�L�*�����Ԫ�w��3N_|R��9?*��+�~̝f�"E��$l��t*�9�y�X�Pg l˔ȵ�$�T����0��<-�|��-"FPm�N7�v�4D�xw��
���a�Z������/.�~Iw�:)�=y����\3��,���\}�R�RlP?��|#�|,=CM9��w�aw���Z2����9��B����+�9g�yӘbfT`�(��Y�)��7��פs�'����ô���y�޲��hk�N"�*8��[TZ�|f��T`ѡ���L����1L�tw��$}.Jϧ�ir �ٝ�MP�jF˃�/ll��?B��F�X�"���@��Cai��(��ۆ��k�_v8�4c�uc(|�E@	o�v�ׄ�@xB}�$��~'6��۞���:�g�V~��kM ��g�w0�o���Rk�ǋ�)��+%̺�?n0�ƕ��.�0rM(J�e��lqv���rc�;,���)�����|Q��S�z��7"�����:J|���R��������<`���za~/ïq�8U�e��G�u���\`ur�H֍�tǡ(��I�k�{J�
����8�GKT�tZx4���ցNM���6W��Mx(c��ɍ����?<����b�lo��$M�&��C)THX�&E<Qm�����|(O��M�t^*�@
�j�î<�޳ҩ,����G`ݑb�X�H���//毱�<9$�+��p
m9�Z/c/m/�5�_y 78�i,M�:
� AOШX��"?m�Z�
�}�
�Χ��J�=)���#W����Uxӝ$���o��$À]�����{��MΈ��)�MEw�揆�I��w��WC(=1�����P��ZζA.���?'x%�4���s�:v�����Ԇ�u��N�}6O�T�7�C1���n#���d7�r�%cV�A$�ۘ�Cm�Nɤ�/�u5�6���?݁��Fh%��ūɄ�&9FH��~0�蠰&���[���?�և��쮷Zث���#g�g�N�j$�7�7��Dɘg#K�c�E9��|�9�Mfԫ-qO!ض~/�z��h��]���\�6	f)��i������[Stt��\K}������e<I�F��T��H+�Xv�F�X���&~��?�г%�G��>U�9b����,�+ rU��2�@�f��}Ȟ`MV�9��Џ����k8�'r����5�~ݬZBj�:�\�Tyˋ{�j���9�nw_y�҄f�ܑ�m���b���ldh<�qw�w:�	)�E1�}��'q��ՠ8
ޔ⡆{�S1�F�0�;vGeڽҠ��~��A;�����d����<��jڵ"��Ӛ��O׫b�v�Q��m���y�y�M�C�t핱N�w�mb7D�Q��kqv)݈8��o�^�Q��Z�L`0��).���T'1�[�p�G��D:X���2���Z�׵��kYS�e���Xu���΃�JΗ0�nj_7 gy���Y��k�l>�����:?�8��L���2�V��Tk���4�d�k����_��*�=�f;�К��������8�4=��r�fe�?/1}�SGA%Åd?�����\��܊(����D��+�Ǚ ̳+N<V�ڞ�P�|\�E��?e����^��q�u�i��]4E�:��QH��{�I���.a��݃u�T�*~aLO�Q����Ɵ�pEuf�v��P!����U2�����zaΞ� uO<9nLG��n���'�^�W�,��$ؿ�u��ȯ&��Y�P#��X�B?h����S�g���( ��V)Rv+��4�-"���D��"I`9\�/^�`wO�)��\+O��DGM�`*�x��El��#���m���(-�}5�|@������ۏ��F��V�������sJ便���^�M�����W������}S*��h�-��N9���>�5`�f4l��b�����H{ �*Z�P�6�&s$J�q�f�n�P9�C7@[ "f�����f;�����<��WghL����Y��(�J�����א���������0F�;��[X0�0@��}"�7��4�N�z��2���,�v8o�k���C��B�ÃT,h�d��0U�*�OC����i�s��/�U�R)[|����Dz�eY�[w)��AE�h"�H��z�Q���!�s��N<bf)�ӯ������xb��U�a
��8.� ���Á�Y5����/����|�V ���?[m\�<	B֢���p)IM�}	������� L��V���2�(Cô�����!�P=�Yx����Ca]X�$�9�`�؇�PN��*������p?�I�m�v����K���=�t�1�C���=�0Y��R�_�p��?�[о=BMҕ��$̌�no�.2�}u�LFD�n�6<���b'��&��uy~,�g"�Я%z�PD�P���W_�X澷	w�,M��j�~/IT���G�>���w�L?�.� }4m�:�!�cߨ�l��j�JkFd�bϠ�]�[Z/`]�i�+3�2o�x����
f��3�tiR'U0F�*V�oF�!IcTb���v|��"�d�����!�7βMm{n_�y��L�`9Uڑ�@�O%=����&�b�((_���a:Z�U��^/?O4^yx�q�(~[��Z����j	O�0÷��'"��
k�}AV�����HB|֪�EM���"E!2�X����$��r��Bc�FOb�j.D��R�t����D�_��D���X2�4)nZ���'Z�X�,�S���5T�`2��򃓺W��!���4
6#�C�h�!~z����-r���)�ɯ���5���2G�r�98�o�Ra���0��]�,J��xQT��� ���7�J"�h���d���V�y�S�r]�A<]M>�u�1�,HΘ=�Fh�e�W܌��7�����v� Ո�@����Q�kKE&���ve����y��4'%�}�#Żl��H�i�����s�_DP{���ϫ$ٖn���F�J*�.8d�H��gr�M(��$@IP��o��rt�Պ�p`|36-g���'Do��	��wC��3�~�2�4������;[��"����Ţۆ��G�O��=k"�U��?U3C�QT�9N��C�M��Ń�/�Ƒr�H��1%�G��b��;��d��Wk�s�ʒ��������^���;�ݴ*��3�
!����N����e����c��o�g'#�ӺS��X2�}=Բ����<�8u�p�eK����m`-s��u������hMdA%K*�ҟ��h��[�UҮ!A\9{*��K��n�q�	E�����a0*��2�0�||[�M���pC7ӱbu��C��X���@U�<�����t��>Gy�	i
k��y:eA�нm�����Ȣ����(<��<�*?F ����i�UbK��g@1ՏAq���э_}0��}��I7r��X�xH�e|�η L�ti��9����RZ�h]���>�2���p�Z6Y����41@xM�e��|�/p�S�`D�'5R��yr�҈��o+-:�⽭�|w���/R�E����j���h�j�	�ƕ�Y]Bt��!��}u�Ty]�A���M1z��P׽��GB�3Y��:�7_��v���'d<,�POU��k���
Q�Ӂ������f�'���*;ŵ��  ���]������ҰpX�>� q��1 V���iW��M@����T�*�.��;a{�y	84+�4� O[�_E.g��OL��G�f3�5���g"�f�BN|7�.;��PG����Y�/�к��OrH�I_�����"'���y���C��{�,X�W�>�u{{�9Щ�/wW]r�P;ݭU�!>@*�y��1b�o� � B���ǠXB(`]$mz���"̗�n��Z��U^���U�:�&W��X��s�D������ZҀ�&���1J(��n/	�����6�Mǔ��
�G�Yk�4�RKEyr4:� 3f�XpC�}��sɧ�g$����WI#�}�k���F�y��· �zɫ�������i�5O�ɶi�-�$M�{�0)�o��}`đ.F�^�����žl�Z�O[A�8��F���*�<9�a�īk�겠�k8�y���*��S�[�"
��o,g�7�J�ط��,(�*�ߚ�u�qw9��2�8�}��r��=�o8���M��,������o�s����ѕ������-��!2;�ƶ��*h��?���Ҋ醍�����R�
zU�#�fc<�v��]��ƙ{���}��f��ȇ�X�����Q�7b�2��Mҋ�1pLuV�f�O�O����S �SB/K�" 1&x#�G�D[O�Q�O{�.'=����|琲헶QF�h��g
���\��]�s!�%�9��UzK)yB\�ol�s���0��,�E���D$�aH���۞����[��\XΫ�|�ݖW�.�:b�g�P����xM�V�G�ϖW!y�(���G����3��e��E*ܰW�2������Ң퀼ůL�!���~Ӛcz UݼX�[H%���0�@f�	ۧi�!v���A"�q��@�3��ۡ�ex"0��ch�bj��}M�.J�<�$���FF��.��)S�Qv1��.1*NC��LE�3�r��������u��S���������"M��S�؄�!՛%��-�\����7UT�Yc�8 xi :�J��(d���@�x�]�zi�#X�K"�k�Q@��Lg�������!\k���1���>l9�"���B�2�]3k3Q�x\� �*��B���C�?��LF���+k�ds�4	��#�-�I�T�#�i�[F1mn��K0��*���sۑ�����h�'��^��k�WfR�9�0�ɨ6-�
���i����UcP���ŧ䠜)��k1��*@+��}����ܽ���2TK�[a��@C:�HS9(�e?�/a_Lj��^�����P��/�kr������j�s6G|�,(O�y`�?bqU�� �|ü�b�FM8f�K��wH��<sJt%�Hj��;�A�������Ik+=� c���\�s�o�]�.݅�ӊ�ݧ�����%n��T���b>"������د�@-��_�E�C4�9W����?�M� ~(��Dp"R��������|��X���p�L.��J�w �S�a��Bʴ���p�x	Ɖ�����2?��I���ܞ��5#I~���@�A*�D�%��H��ܸ�ܘ���K�mϿ�K�8	D�2�(�2�����������'Jɾ�.Z��Xe4�Ķ����T�M�d���@}��ʒ�\QU	#M�w� �ʜ����a �6��t�-L��ߖ����!;=��Wv���Vl����������X��w�֪����P�����b�����6�.eî4w��X����&�+9Ƞ!��P'Ck}�g8v��`>�B���:T]��M�O<G;F+%��6N�4�����]wg�H�c|-�c��dĨ�G��f^�RI�ozs��a�r0�O=jb�톄�j��J�MP��� ܡx����͑8AJF�6����?�0&`,������������☦`U��ϫ��-S�>��ҌR���6sj�Dɚ�@l���p��;�Ҭ��90p���4�����<U����W3�5���TF��@-�%ꦓY�|��S*�1�]·��W⵼y^]m\��Т6�T��KC��T�El��j�v�"ujX�d����	~^�֥��I�8?���N�1t ^�-�f������Xq�I��쿵�E�*�2�4���x:&|�J]���g���d��FwJ$sG�q)R�#��5�3�pb#�#9�]��4v
4�>u��6/q
��9ۧBŮW��*Ch�T����N��sИ��+�l����@��$k�*,{G*9�|ef,���I�X!o����:�B;�9r��l�/j�����3��Fq�D���ֈ#q�T9�%�2ȸ:�9<�s&	*+��*Me���(X[�M��S*��E��Yu<ш�cXE����w!�f�;u�`S��X����(�wV���3�{=|t�8��i�K�#�J�)����,�(r��9|7=R!��lڋ 6���R2��}��P�,���Xռ�v,�07���������li�$��ғf8��Aym�X,��ƙ�6�����	���ґHl)�;�ǡ�Z楗�Ljzd�9T{&�c�f32���يs��e�b����5���i�P����f�y�СKT��$'�Op�ss�y�t��s��X�Gx���0���"&�&��)p\C=�`�~�#U�]�l�r72�4&Ø��b�_;|�#R����)A��"8%���M�Ug�^��}�G���ѠF2:w�gq�eq�P�Z��]'�sc�|�C�L�$�;�s��H�H)�_��.f!���W�b7��"�K˖*�&6k-���R'��dPw+�YX�����m��z����iS+@t+C"��c}7m��DV�Q��~*R��޽K:��)ʖ�	 4�=t���e��CMV(�i6����"�N�W�	4��!����vHR46��� �0�����qNs9��-�)�� �@����v��'�O��!���(/�d`a#&O�B�|�lȝ���_�>>�$h��G�7�)����'A&H�v���%�qQI��>�I!D�`�ͳs��k�$��,/o�-J Q���`��C.XX�o�t
��M�c ��X����l^� 2E:�}�Y�����Fؠ��L���|y ��L�ge]��m⧁����Q��j�B;-w�`ϩA�&:g_��l0n�R�尵"̡-.��W3"�:W4�<����T�;����О��͓��;S5SIKT���b�Ǫq	Ҷ�L
핖�gz�t2����^˰��m�7�}8s�e:�c�N��Y�!>)�H�#�XW�zR��6�A��W2��b`���.��.	��\��.c�~nN��\I@Om`��v����4S�vp���-%�K��EJ�p�	����2����}������D+�F�Z��&����S�� �m/R�зF�k%�����8��ߦ����� `���A�m����Bn�fp��;�O�w�$8��JN�o�����89N�)��|i��F��æ�@�� /�+��E�����XL���Az#:�o~P�BÐS�5@�"ʫ<zkХ��u�Di�k�Ȋq��������a��2X	��pp���:,���k>0#܁�%p�-��2�}Qغ�a���	���ٴ��R�`��3�8� � [� ��.��0L��7�BBj�r�����!O�����!��Sbt��v`b3��<_�D��+1Ŗ�8g��8��ǳ���r�>3����1�i�=�@��F�
�Lé�F"�U-rɣd�KB	s�Z��?	Zj�p��Q����Q���}�\�V��T
]���i�J#�>�G)����!i�#��>��3�
5��Y��@�挂��S,��G�wd���%=�6�>��#E�(�Bg^Ԑ��j�����QUW�hX�1�t=K�UQǇ,#��N�N����;���<�/������AN��U��>�x���4WrF�����q�գ�c"]z��+� @���44�'�p��C�Z~�]�Hi�2\�T)�0@�L��GZ�t��-�_O����xG��:5]m|�<�+�ܘ�����Ȉ��O�Ɍ�Q�/�|ɫ���h�+�J��?���	-�S�oZqd��␴U�hP�ӝ�c�9d����.�N����`���vK�a�;�ăs5�o�n�湿pT���t�L��_|�����o����fEeXhZ@�N�}q��VZ;�ڏ��6��w$��q�6�Α��.̏" �]+��W��v(�����黀" �3�Q嵖�æ��V�'c�Qa�
��^�f��r��1��Օ�y�]/@4%rd�7B/��&R�|r�i�$e	��@�����NcA:��T<P8�)�,2R�=�b�s����(���<Z�w*�5�j�ĸ�"�~�y����$���Y]Z���� �b�zۂ4n�	*�	�M ���,rZű�K� ęF�-��Ee`0�8��<�7���(9�4-%'[�>�\�����8q���S�,i���>��f#�}�#��*�|K�u ���,�^�f%<��il���T��?Q�`����xL^)[r�Np����4��pϋn����KVf
������c'e�1$.��� nP�O\Q�D�dS��w������A�4q�H����s�H�{I��#�Bf:�#HP���C���	S���z��r���%N(�6h�W��A��+^yB2O��g���|#Ҵ3�/����ط��F�|�����2�==�t�]�2���x�����nCl��S�e�.����ǭ"@^�Dc�.I��^[�Ӑ
;̈��6@9rOs�$#������@p�i��n���s�g�g�HeM�Ϭ��츄]`~��d�@5dQ��5J\���4�}Ek�� ��S��K�j���c�a��-^�e��jH3Hi��5Qs�f�kW� �/اm��j�xZ��mn��Vws���iS U�͜�p�R�����J1�̙u�P&���g8�H�0�ߦ]8��EF�����rMh ��Z�k�W7Bm[r%�/*WBs"w1�V�e��,��5Z��9���`sOy���i �߁N����*�D�$ݛ��� ���[��j`�g2�*�e�q~t��N!���_���:-�m�^�uQ��r��*�I3���R)�9L�m�������i~E�:2���Se��H�as�s}.���5�Q&�$����������[N����QI�(Tn��]e���c�8�o��39%ƫ�,=�i��,����d�1�j=�L�I��M�^�MR)�]غ`�)?��[;i�`} j<0��Uh������QwA�$䞫ԟ2�-'��:���QҤc�ֈ�q�>����B�Rc�T��)��49�ʰJ���ͥ�D����������4�����$�#���1 �sBeL�y`ɧ�������ʓ�T��PZ�#�O]ܥl`�M�y4k�[1#�?i�ڟF�vL��<�\X��$q�K0LGHč{�gP�8��_'��*��U�����$dlqJGФ�\u�u�ۖ��UP!h1u�����@���*�5=K����[�	�&�&��ck��s),τ�e>�������:�h
�.W�Q�f�����Ef����/TQ�Ӏo��&]s�="�o�B3��r��S �.?���Vl�Hm$�vZ�����P��q�}7zia��6�C P��r��>[�r���`%��q\�L� 3�ɏe^QF�����}����o+����©���K8��'�aR���9�8��a���9�r6��v���C^!D�U�6
��6�r��@7�v����1�h�ࠃ����ˋ�^� ^�|o�z��wɵJ�ǽ�y��4#�ZjB|#<H�i �]._��,`�컺��[�z��Ecs̤����@qo:�ϰ�1"��qlEb4�Vɜ���*�|h���k,XהP퐍O�ВOË�	�xnIs�?u�^[���B<�8�m��\p'���`:(]�B"IBE�;c)G�ж)_�m$��Sә�Fj��a�`��������~	�?XZ�ʍ�T�2�'��8Qd��z_��,y@���[s(�1z�~/4��_��o��M�.��,"�$�:r�b�*^c�-�UT��yr:�U�	�����۱!YY#� 8j����:���!��+Sޑ1 �Uj����(�ލ�b��ߏ
���U_���.�����E��B���t�:q)�54�ʭ\q�D��j|^�1i	攋u	����n�@�l�����؎�]7�s2�mS��9��?���$��fi\A�����~��NQ1Nb?�+F��yS������4�|&���g�g����U3���V��/�Ƣ?u�褺5�xqѣA�HX6e�AS�X��HK�^�ט\j��}&~18��V$R���f�N�X�KJ4�L�1����%h�+�,�[=4������b�����j,	A�-X#.M�W���s��0oN1�ḥ�>�����@��$#��

,��b�9Z���`�ذ��`l���<4��±��oӠn�ǈ�R,ޙI�f��+{��=��`j�`k�|[����lMV�@#G*�$S1��E�~�Gi�o�5���1��d$�����U�4��bb���w��g��śKV|���P$�ca�wې9N��4\��zqA��[�.�\��A,D` `_ۜjÈ�;�73�C�q-!1�%��x�l�ς��d�~��$Ӝ.(�D�$�Z��q}WVvy�����s�!AْR�?K7kx^�w�I J��m�A�F8�K\6�^F7�P�V�th��{��K�@miQ��)���b���S�	tWij��tvfQ)�]�fM�/ݹ*x�-%��L��Z�L����0�sv@����V4�#��M�Un\^!d�ߘhU�oX�:a(o��3z��r����E�D+��4]��a �08��s�8ZS�[����l՚ir�Q�5�VM�L�*<�2r������}#�`)U4f�]�C8�B�Ü�G��i�@�܏FkX�@�� ��i����2�1m�kY-+�@�)��؊jX���yB��P�r%<nR�'[C�h!6��*�^�Y�L��2l�eS��z���/�1.�[���__��?��͛۳�IN@N���r�KV9'#��|�>3��ȆtG�LS���<X^m��ۀ�m$Hvd*�M���ؙ�E���-i��ן6K�!��/�8'/6P�0��o��ͫ-;s+����\�>xE�sl��j���n�/VK����2���%��*_��`Y�����_��٪j�@�3���w6�ږ
i��E��G1���|2�<��.�ɇ��?�Hm��P�c�3�/���"'�)� �U�oO���-Ϋ������?9�����]u�	6�+���L�5����� vD�P�CRy%`�qa�|�;��o�g>�h3M͒N(U���֍N�������U����6i�@���Ksc�+�>|0�4Mοg�t#?�j�K��[�?e��T����=d��{bƬ�}�X���L��G$�Q�|a��(%�]K�֘�7�bȡ�O3N��������6�(N��J Q�� ���r���a��D���J�p�AFן�����xa�\�i�3ÇѢS|��"���Ჾ�����oEau�$%BTd�S!��s�{v���X����Fn��`S�ٷ杔��}�G8��3EH1�WS�AG�����m�_����%�͉�SHj���)��l�]O���N%��s�Nyn�TN� *���;6�O�6�� ���(��vC��A�%B �lN�f�M�{W�u����3cՇ�P�}T�"�%��̋5��`�mf�[���
&��E�`4'�H}h�����T��[���7�9歀��7�|AB��zP*�:`�^2�����_�����q��f���X����o���9 I�*T	+�=5jy�f���Iߜ��MT��������z*�7����s�U��/4���F<��L)���,9��5�����W�k~��_���e먏�l��8�j�;�ҷ�k*�.��w�F۞+[oTzp�U�/��?I�%;�
��6ʭR-�k����������k�v��8���w��>���r�2�ܗ��*,*�Xh�4A��_}���
4�f���[Ux�c��0]��
�O���0К��.������t���+����E6a�՞����k�T��j
8*2"���G�`4�~��o��iH��$!)��0gW"v��ce{k��C.���\",g���51��)�;P23n���Sbol'E̮�M�#xrN�`�Ⱦ��:�'9��`W�T��]5ؒ� ~Y
�j�\B�qZ��[�N�aR�<|�&��J���"���a~<�byJ�2�t�PG�V_f`0���qWa�]���R&�R�"��Sf`ش��1���A���j}���4��hG��>%��D�p�����ȅ�_#Π��L��n1�_��a�W��͵#^�a%+�Ȱ�])6����u�"K�������yņ#_���9"d�*������89f���j�����⌁$������m�7��և�������b���s^���lI~��"���]d?;�ֻo�-1u����"o�?zm�f�������xs	h�g�N/L��&�ߧ4}�ɴk��))��>��9/ŠȨɪ�}#e���{=�4�ޙ�Z��$댘j�R�i?\�d��M�ƏJ�o,玃7�6լ4E��s�q����Q����\"P�2g��^��{��,r�u~���4<A��&l��B���5M0�z��x�ʦ2>�&[���)W�;F�����jN���W�
j�2S��#p"�q����� 5K���Zz��]���!{K�l��A����?���Q}�X���G��L��![��v~��v� ��-�t]��\e�*J�	��L����P��F�ʓЩ��
�Yd�̑R���(��������*���̰qs���0�;��k�+7��!�� -�i�("C.p��4�M{;r�A<l$��t��B�˲[ݍ��\A�,�W�BPq2�-�qA}&���WO�xq����L�:H~t��W�e�n>�>�.�������wwdl���RL���/��7,�ݳ.�D���* ���� >��V�1b�ě�$C%X&;m���B$���򏧭ϸD�Y�q.�O��6<�%�V�df��]KB���ߞ�y-��މ:m�7"���"�Q�d�=�̕��~8��`ۣ-q�7B'(��j7e��~��1u��v9��Q�37������6�n�J��w��rpH���|�!K"� H�t�$��ZpB��ȼ"˷D�}��[��i�ԗ���m����ݖ��T�$�E�Т���Y&�>�Ð�ԩ[-��Ysې.�g��^�}Cd@F��g�Sܥ
@^��7��SQ߯�����mշ�-��4��֬��]�%+E����0�90� �� Yw��t%�k;8�14[*�^������[�-��FX,�FK\?U���L�f��:��?m|��%�-�K~�*���3�aU�
���Ǐ5�/������M/fR�.�p��ar_�F�sT[d���A��7>Q'�Y�^�)t1g�ǖB|��\�����RXT|o�%��� 	�`D{�� ٰ�=ܢ6Nc0]��w�ԛ/!�N�eo@Z�Zu�z\��
»¹`叄b���[��/,뿴����:W$��sj�=Cj�I����:��]�����gz�N�{ʋ巌��QqYu(�A�Qi�'���g�T�!�ɞB�;-ڍ~M.�{��X ���� Ы�
��|�Əb��9�`����L�F���͎6;�6�U��Z����
�x�x�J+\�|S�<~�+i�z�QoW������R%��?x��I���#D�QE^����\,���#���IzȧM�MՐ�Ȼ(WR�����I�E��	�i�`�a�mٻ��rv�@'�7�K�_����@V�T���j�s-3w't��ODE��f20Z��@��R�d�*@�m����u1��bdnHM{i$��YU<��^_�2�H��+�~ǀf�w���S�������4�'�eO��Q3z�=��}<���l$�W�N�P����5�&ޥ�ur"���V�ROGS;ʴv(���<��`�vjE/�5����� N,E���:Խ��p �H�j�����o �|��2ES�8���Z��. �e��w��d�m�-"�4G#� q��Y/�wNЁ�Y�(�B�>�u*H���I.�]#��u���:�n���{�Ǥ��y���5�cg�͍�I��zc�V�����bv�w���@��
(Ift��z����1N\ E]���!sBݯ>�i�(��2�F	2>���;��U2�����JZ�]�tZ���E4��O�	��x�;��r-��>섷�?7,��J��xi�V޼ŗ�l]Ŏr:aP&��N�Q���@�FL�l��`���B�Z�)��������C�D%@�i�M�;��zn�Cc�a�� y���*��	H2ͽ��Փ�>J�ɉ��\��sǸ,�i.Sq2��L7�	:k���ӨGj�#=�t��k�
V���� 2��I��S4�O��o}�p��u��/��wo�6����QDSj B��b�Dߵ�!�%�d	�&V���*��H���>5�1��b�@��̖��^���
�q�kb��@����+ד�h6祀���'{<�վ6��&�^�K��h�4v��1J��REm@�Ү�l��N�l�]��8�\�cr��Gar,^�gy�>u��u�
���`��m+�ڦ-�;��?��PL�xzd/�mn�ia�[��z|�������-#%�rۯ�z,�0��w�디�T@��㡦Ad�@����xkK�d�FU���b�RFR?���NP��A�!�;'_9,ו�L	�13�f�nu�s��֙��M��m��%�ߘ|H�m*�g�&x.P���E��F�c��iα�
)
���~1��ɥ����B0�����9�pnefq����zaP��s�����<=w]:(�y��Rc�\���c����i�t�R�(�D7j92����dt�)+
+��;���R~�f���ʫ}n������-�n���h��.������o�%��L�SG'�g�����eZ���(�-���1v�4Vz�\l����t8ev�2���L�M�A�p�^���,Z��7�p��\�L�=�f�Xs!qd��n��7M�eSvsNػ���Md��+�_��(R��{����d�d&��4k������.��1G�`NU�z��<���UY��8�̀��uJݨ
�����l��2Ȳ�5��(��5��g7��u��~�S�Nɵ�(��W�o�+�yO1h�T6a�վٰ�ŘO�ɊB	�l��� 
��~v�6�~)����̣�B\p��:u�w�vPr�	�i���Ph�ӟh֒q���%�c��2�j�'Y~��%�y&�$�p4<�/~ڃ4?T�|�s$et���"]RyO;j�������{��k�#ם�D���-.�O�Vv$T��Cd7�M
(
���i�ս&��Z����)^��e��}�@�
s��[�z4t(�z�"%�������� 	m��p`1��C�xq����n3bգ�OM31C0��ZhҎ�Xv�^H���x��~�	�W!���d����2��檊�h�8_Q'��_������M��,��A<l� z����R��Ate��PT� �~<��g��B�&�6����Z?c������9����-�n!$m��t���S_Ks�P��AB*?�F?�tG�rV6���T �ؚ�"�̡ğ��.,WK���<C�w����0�.}y����=mF����ǂ�m�&#r��w!�H��Ѹ>��|�%�=�/#Iu_��p'1��v��r��ﴄ�[Nl2$����W��&.{�x�1�~h��u��]F�\d�]I?ʇQP�˧����@ �Y���i�|>��zȢ��K���4�f���<�3b�z��q���z��:ɨ2O�bA���j�����li%�DK��5�5�H�Z/�ω3��a��G��>V��%���Lf:�%�t��FsЃ`��c��'�EL�a�7��@0�K3��v��0����
�z9#���V���0bлi��]{{���E����ؼ�6~���ic]0 �
�f���/a.���:V��j�C?��6=.���֋�� ��M��'�X�G��f09�p��#jر[�=�����-����sd0�B� 54[��A9u� k;��b��n���v�^�U廍�D�B��S��Y������?����5]fO�F��aカ�Ҋ���}�;<qt�D,Q ���;�CJ8���!��{܆{<x����cU�����8��Ә��]�l?�,�m���Y��`r<q�~�������r��J%��5d�9�c����~���`9�(�����^�T�ȫ�xo�����zc�����;F1�U��*+��ჱ�S���m� ���;�O�u"=�ԡn�6[%���ZZ[��K����n�>+�0��t����1�YH@`\��?��M�/9fD�"����$���������V&���������HZߛU���vs�\.@E�Ȃw��}g:�f���G�d� �������w^�݉ǤOf�W����N�t�uw+͝y���_zq�A%��O�y��\�P<�mA*q�Dzu̸��D~ia0�B���ċZs���<흯ڪ� '��6Ʀ�]`� :�LI�����mf��rX@M8�Ə53� a��Y���?6�4h<��J���(~Mp�lj#�D7d�wA%����x5;K�:2~�	�4[~h��j$��0�4�0�&L�ג���T"˖�
����` �����p�z���e���F�m� EO����Ql� �cP��Ľ�zF���z��;��h�M"@p�V4j�݊�G����RP�p��K\m�8�zFj���Hw�&�e��F�#h[}绯���e���j��n�I��~��������l{*a���յV�xz�"������Z��"i��cF�?����x��۶U��x�Yݞ I��XjN�9��>Dnq��|��R.��a�C�ҏ�$]��cn��"�Yŕu96\�W$!�G���s�	4(*��zr��h䙯
V%k|�T��=W'�I�}�JZG�q��nM�;۵I��VJs0�!�{������e%�/F�
��N6���JV�&�Q�	� ���1������� �3!��(}�U�/**C�����|���WR�F�Оb�
B�v�G���?ÝOY!N��ą��wZ�NL�[��2�%Rz�fn�c�;?��2v�"a��쐓�+HR�]������69s��so�Vi�Q��A3?j�BX�u�v��s��f���ylBjEMG�J*��R�aβ��?@��w����P��;4��SN�'}�"4/Y������U�½�T�gn)�c� t"��&n��3���0^%%����WL��P�����N��|�:��������� $?Y'�x�bڱ���$�z1Z�+.Znta��������A�0Gd ��B5���7J�{��%5���m*)OaR��$6�3�� T�`%�lY�p!�ف3��:4��SA�z�L���� �<6�N0A�����IGZ��r���ҫx_=؀�>���.��oXqR�[��=�m�U����2���D��X&�,�ʒ?��^������1�]�gK�
KL�QbS��E�@bK��N��f�3a���E�Qڊ&l2S��_v�Fu�w۠�n��I:7Ò8ZW����,yuAY��i�	cS�<#`���D'%e`�%����s��Zy�=�k9C%H\ԑ�����}��ņVT���C�ˌ���ݔyɸ�n�!"ב޺cK�=�Yʊ�Y�ūͨ�>q+�g\_ߢ��O��������a���8�)�7���b]6íY<����ON:�iL��u&��F4��!@M��p7G�m�ҏf��C
�y�鼬���x�RU<C�6�!�W3w����b&�X��8�PH���"����~�A���)�G�{��ҹ�-��l�Hc�$����|�q/�~�OI�Ũ��G!Y�V,�x��?�03��y���M��G(ޙP��� �ɠY{��gDw;X�I%(�� ���	,� �� �D�'���n�"~�����/G%�L�3`�!R���;�A�u��{V��E���(z��B�����;{��������#���f`��5�q�D��Q���kl2Bxټ��l�i��l���.��X�[4����J�~I@�&ڳ��U��=]��#	λ����t~�ҏ��h��tx*S�����6���@|�	pB�a����~�`OƄFn�e�QvAPo��5)�е*U=��e�wt��2��办I��/A��8)pԺ[LkL.I����?~X��Lk� `P��/+6�����*�o_=UZ�;�4@�:`�0�G�wf5�����r �I��j�-�mPx˷�/��Z���E��Ӟ��H��v��
5#�h.[��P��4d�M%/C�rK+�o$M�Ϭ�;�Dd�%	�P$E��}ׇ�����\;�m�=GP횓E�X�QΫ��K������-�}��1"Rj�C�� 0�{ ��S2�fy��\A�Ϯ(��եÜ�߂�m1�wC�\�^�-2JUwx���=T6��U����^gѡT�������ze��!�.�Q����l�i�5��ҡ��'�߿w PLwn��80\�� c�^�o�g*��W~��a�U�hF�*#�|_���
�ޮV@���Ῐ���/R_%Q�m~��g���Ub��!�PI��<�3��V�M�k%Ց��Wѕ�	%�ΘZ������(���[e��^R�_N��h����z��34D�V1͂�b�E�*�/;#��z5[�:���J>3e�A�K�.z�}���!�9XX�WT�
���͐VЅFB��p�3����:�Z��d�Ц@t#�Q%��	Zfp&e�*�9��r'W��̦�ž,;i��15������;p9vvƜ��r�e�@i���Q��`�+t�K`�)�½U`H�f����t�T���*�3���D�z[��mu��� ���J�����La���.#L ��/���p*��E�G?�s�E3��T���{��H.�,�+�Jw�G�0�3}���yjG�f�����C��<�-P�Y��!����m�Z�Ey�H���Yq"��ϭq���
q��v��A}A��<{�ǁu�۫��5�.�[f2z�]\�?0�?��9���5 �6�}�����Ơ��\i����VB,�W�4?h�?�K��¬-�q=0ڴ�{(�y���H��7:N�t24�?���w�&)�s%wU�{���
%tSz����D/����_VP�I��s�B���z�i�'���~�"��7E�G螌�ry}���O���u��X^g����m�IOq�������9STlN�n&4�Q�FSZ��0Q���Vio"cu���=����Yc3p��"����Ċ ��}�ge�x��ya,�1�Ïh#`���lۂ띲�-k"�@�n8p[U�]!����[}�c���P&d�KW6O�iF�w�E��"��\�p��wd?t j&!�7�G�<]��)��ǔ��#�쳅M -�/c��ǨŲ�Ȑ��+E�r5� �pxK8���p�����z��Z�a=�D�a����TU5��p���8�����г��T���ܱ��%��;ݲ}M��h�xĪ ��q�`f뱽��l�)�a�o{�x&$H�:3A5���oZY �=a������b�ڡ�a��%e��B����+Qœ��W�b87�m߁����N�v�Y��z��_`���\R��y�.SX5�̢��L��M���Zk�=��@�A���y/�'���ЧB<^J3!�#�������n�Y�v����d���ś:yDW��?�y�(�yy�bgIH�r=��"�8��Y�%�P\�<�%���;+Q�2RT�kq�$/󼑮n�7�DԱ�M<AҎ���麄F@�ư�B7���q�t�?�R=��%/E}%��l�C5�na����<[Y�
C������X'����K�4U��<!�@��	I����KƦ��	0$���S<RPZ�:��]�G�����f�j����:Ɯ���N��<2���n�Hr��D�Y�g}��	��#W��Us����J\���(�N3���d��MM�8�AG�5J]k��o����ߋ�����rH�����vQQ����4�a��{�`�q���a��f� h*�m���}*m��p��C��E���v��ȷ�,Y�M��?=]k-�ۦ<W��b�m� 7Q^�iaN�ME]�9���ۅWS���D�q�:l��]\��"�q�a|�O�:P��
��[^�\�Te0�!\�&�M�U�4Ȩk��0���9�oL����lnL7��
�
�����r%a���NC�T�U{�9�H%W"ө�����[l=�l�����txш{�^�RB� ���Ө �M�v&���e[���G�jzO���-:�|�H�h;�~٥���j�W�_�%���o��l`t6�!�����9q�_W���:�ſ�7FOӮ���M)�r�k*r4u��{���I��������~W/�)����������e�"���I��#I�_��t=��ʁ�ٌ�0�i�|)���䕏*5�����K���*��C���$�0��2S�	�bCu�;O+�L�V(e�Bm�P���(ܹ�Vy������;�����66��6��@�
� �W�^��Y�����Gп�U9�P9�ȩ&"f-���}�K��/M�C/5������<�R�'Q�I���,䄸��}��̈*M4e�NJ;�sv���X���ϒ�d
�3,��zn����L�n�G*Q���Qsm�^R�2"L�;5�L'�<�Mْ{(�_��m��3$����|�V����0�#�V��v��
@˜�N4dN�a�4��@����ϻ�v���8�,��玞�@�s�!�e�w�3��\贮}ڗ%	R�S6"�<M.��ɺ������g�>��� 1Cd�Z�ԇ¤�l�)ﯩ<Z���3��j3����y�º�͝uH��7�ذ3�hM+���}"�|NŮx�&I(=]��-L��-�V ��D�sN��d��;��������_���j�9�~ *���V߄�/�C��8gZrS���y	��}������`+��Hm�).���i?�z��;�2�I[�d�Vm/k��&�W�K��vG�W�+�+�b���~�G]��*A�f7
3��K��}��F�]娫��0�Y#O$��Bs`4O2����������	�4����������ZF�l�Zx�O�8]MA�S��C��N�om�}��� ���-rk��E��P~�ޡ��0p"�e1�nmHμ����zF�o��z�����<���i��ل$��ک�A��d^@J4��ۚ�m�-��5-����YpK�]�l��B�T�n�8<~�p.�-�H�_; k�>9F9�Bt����,�0�2:�?��BW��QR͋.��)ٞ⪲
�I���{���Qc����P�1Z�]{d��h$6�I����h�}$_�ʎu�d��L)��Qw�-��r��U�$�A����ɸ�[p�������>��
0F0���E��9����6!��~�Ƥ 2�*K��a7c�=�߉CM�?�5ͤ۾z�*�lz��o�f�0��w_�i����Q��2����/�E[УU�^gz�q2��H�xY��2��7��}��|{�VHO0��S�27�H;�d�\��TI�K�`ڷh�_�HEt���Rj5��
V2{��R����楹fR��`&��7��D^J~r�<�"Vg3�)\��^�;Ӣ�6���&7�9$%���Op�&x.8�N~��}������_W��?~�p9�L����\� �hj:�&�E6��'$����a�,�ܟ�?���}-~�P�-�B` ������Z���}��*�v1U�q�0�5ߡ8YOb#�=A���Pr�BZ�@!����+ORʐr���c�8���[&TE0?�-�l�6���U���Ba��������tχ�b4�xj8S�;��Ч)�<_L}��׼�Il3n�~y���C�T���>��e�$2�'��Ɲ� y�� �,t|GPq\�gՓ�,�s[�V�E���DO��$]���O`�`�}�zR�_ߙf��Q��C���i�<���4�Ƿ�O}v�0�bT��[��ul}\�-�ȕ2 �,�]���Qq�#�'��ѼdWu��!M�j��:b�sl���k��>ݻ�'�nȷ��xp�%�_~��?����jH��fjtQȃ�ޡ���4���1�������}�R��7��\&C'��B���L�{mw\m��ܟ9�˰H�,��k�^�����nhS~��_iH������[�-Fs5��{��������1��4"���7�?�D!�C���s��(�Q�Q�_�x�rTs`ÕZ?�rL����簱x�m1�ՆP?j�/v�8��/*\���z�׭�T�<�(G/����P|b*� ���"��i��IVM̻�8H��DE�)��m7{¥�Q�+�b�ۂ����<��ׅ8+e���Xo{���Iy�\zW൳��� b�7
��H������ˌ�Z(�s�:�$9�Xg����/F~���g{�ȋ�/��-�%�l��]�-Jq�[����U��,�}���!��/�w?�m*nB'`7��wgp?�A�w�3�g�]�M���PA�Fie��TI\1�c{,�B� ;�wHY�ӯ�+��Jy1}�:�u������I񚮋	ߍHD^����/�(�+��c���2��.���ZfKUK��tyz���JX�MYz''7�e=7��s��]��1�SB�O�t�a˳��3�R�� a�"Ӈ�6���yj\)�XSW��g�k6�M�='���ւ�f��~%�� +��a�j>�l��L1H��*�pZ|������˷�ꤥ��r���LE�w����_ڼ�pUlr�	�Va�5h�dW��Ǫ�@�f>�@4J�aQs��$c.7�,!��ү��Ҭ)g?s�/��ޖKK�%y]�FN �2�$�$�a\n��ߋ���ʙט��Q���Si���Hnh(	w󂟣X�n��]�����)-�x��h� ����Ԣ�˧"4�0����U�E����:����
hp����Ǧ����"w,��׭I� �Ge5ts�) �|n|	�`+�����<=II[w�X7`�|oQ�T���m��M��:o3v��I�f��k
C��|-P�r˗��61?��<��K2E^�dCm�p3������>�C�G�V��Q��.I���6��)GN}�b��.��0�|ɊŶ���߂�OO���1��x{�3�`2���ۀ���%K�2kb����Rz	�ei��}3I���G�?Q�+��	�:1V�;�b��{�(�\2^ٽ���# �yO�V\�U��D2ά��T����Vp�j�?��ڄm
�@�C~��կ��Ț>sgqAW�5.B>Uq��e�M��C��	Y�[Cv�j�I��ȹ���)���U��X�g(Ԗ�F�@$��?0�а����?�?\@�˦/����u��m�g�K̺�Z�)ρ}�@jg�'�-5�7T����#����F&\�'��9�:��Tf��*��d7��Ϸ�6�NE��e���P���"&���wl�UC�s�m�!�%��y�t�P�efA��!�	$�Y
;�`���8K���Ѹ����7��(��73�;�#�x�+_-�yk�.�յ�Lc����tf`�D�]U#�iC��OT�/�݁�����C�i���y�LH�IkM&�ȶ^C]=��: :����Z�s��Vh�F���5< �Ĕ3"�U�jrI&�uIh;�x�6���t8�m�f'+���՝O)O�ݢ�LP�jm���\<����![G�F��p��� 1쟏p1nm����;�ω1z���-�;Voo���뀀����k|ë~1�a�˥��� T��X07�"��]�\Y�2:k�t�K�vk��B�n���G�w�[rW��v��S���}Ol�6��ќ1\��)��>|Ib��6�*~��1^r@�4���g= ��0��- T�%B������?>�(H��Lބ��JBiF�[��x��V�
r�P����%<�9��uM��kS��*��$���-!&r>w(P�z�A��D|�z�����{�5�0T�7���^D{@Ȋ�N�P��cB30���ޞXL����/sm$w�� ��k��-b0t"�C��W�����92��l��<���c���.�ޅ��~�W?�X��@��KÁ��"i�||��{q#�91��m?��3n>,0�s��o-2���h " v�0��{��A�y��M�3�\�2ə������u����Je��$0>����<���^E��[`�J�m��e�"B�+��Q�X%bs������+�e#��ɚ`i(��"��>�&�X�[�H�a7ű��P�ȅ�ͪ�>��������R����ڪ�h�=g�4?Z�d�AZ0p(8�z �u����ж�2h�I2�$4"{t��?}�Y�q7�"�q^/����wǪ|���Ԗ�1�U=_��>b���ރ������˴�8`�!s)hޛ,��)�Ԙ�����7Ng�*�tlК����:k��C.�Wܽ;[׸�zIC�2pTw���M>`���k���3�_P���RȻ��˚��(n�R�:m^�۱�ťa�9α�����4
���YG�KbV/�E��H�FFnXܭ)���%o��T�Y� ��V_���(F�L��w2��U��+��ۄTW�/A��V�_i�(��S�}�9�b'�OF-�A�𶥿��2�O$��|���:P�"x��zIw���[ :�O�p�,K���������mRa�(e�o�u���j
��*���b1�B鱰��d��3/,u��`�jP�>��v�z�K��ӫFJnyAV�>�P��ɛ�}_��	mm�D�:����k9�d��~�<�p1h=��i��G�u��/ 0�%�*�EA�B��_$����h�������'����(A�8��'��%�_M�a/&���
b�Jǋ2i;ټ�hj�ݱ��W�y�l���<��3B~�^Y��#T��?=�s��4ko�L���3n[�Z����^)#��@ϻ��Z~������h)Ѫpz�k�Z�v�� ��8D2�O*^'�=X�.3��K�b�I��{뫥z�csw�j��VX,�۩��w U4v���M���?$��F֘��ǲ���3� �Kt�i�8#��iԯvGr��Y��i~���6��c��/�4��6�����n�����'����BU_:�P���a@���3�bo=��^�YG�����Iw��}�
q�(�>�NW ����ۃ��`Gr�>!���ge��2��i����B_�fj�QV��d~�Y���:�e��3�F���5	^��P�w,�`�D5��@�v���$��P�^5c�+��t.�G�C�VN;�JG�$���g��)W�^�����V�28[��34ᵻag�F要�C�w�������9�90���l6�H"��|�@��v���l�c�
xB���"̮�+tnC��y��q�fF�_�����M/y>o�B�
�Q	�XL����qd(�xv��H�T���@�ΒMo��C�y$]q
I��e,z:�R8%趈��r���x�?>zk*=��P�#N'UV�by��Q�V��\<شZu���v^J�m#4��.	Y��~8L��
��P���hW�k8z��g�"�v!Ơ���*�CS��LB��⢸%��C��!Ieـ<a3&[q�*d�ۉT�k��*H���ӄ0q�u�:g��w���PKu���C�p��Kbo[�m]ZVT�:���J:�&���{!Ph �D��Q}�D]$���	d�)񕻗�Ti��v�|�������a�Fu�� �Fƣ�{�T�\�>֤��s�oZM�T`?�\6��`3	l��y�'B:t�Y�(� K��i�e�ur��2�3p�;��5�.�^wNKp=0��2�q'��[��]J��$��hi�j������������`�r����ۍ�^�����g�.��қ�
�����!V<�����ǜ79w�wBXe����`��Z^����:=����#	�`�:�Ȩ�&O��͌'hv��o�]�Zѩ�ǆR���5H��F�ץ���p�������}0O��R��NU5:��k��G�*l]�f�M3��G����I��Xz{l@���f��1F��.�#�хS��;���^�7���L�\P4���|�5
#	�V���KY�9��D7{���ᾑu^�e#�g.-�%�M��Ⱦ3Ԡ��?'��9�3��jLK���Q0x��H��t����
bjg��6�OP�@�z������������t�$�	�0�����B�j�\��#��:� q�XclB%I��1h��r2�j������nRV4{
c��������#BYG��ʱ�ʀ��a7��Y�8>6� ��%v��'p�~��b�<�eݗ��-��+����(��
0&��!��7ƹ,{�i�P�Ix�@���WHL��c7!�?q�:��a��JV��>m��:H���C�§���e��O������Ujq;F�ѻ
h��e�u9�B�U		(XEDJuT��;��[���=�0gD
ѶCҝ�1���{<Ь\[:��ÿ���G��������(���� ^/>gG^��s���U�G�cM��F$6p S|��:�g\�n딟��3��O-�j��8�"XDv0$b�$t�X����9�/�A����(���|���Z��I+�y��RTۆ|�BFD96cޒ�y�C[��D���s�F����V�W���I�,�P�_�����p[bw��M8���,��$*M鲑��kHcG��*�l� L�e��ǝ'�`��r�eq.alP�������CyB�>��/5躅).�WMV����#2��?������?�+i$i�2���3�VH�!|�v,b���b� <���;01�;G� �/ G\���[�N�zg�sG�E!Py��j����D&��b��~��)�<�������-:THʯ���^긢��d���:<٬�z�av��!l.%p(R��@����w�B&��
�����X�G>Aq�<�ث�lš�f�(B4�4�ER����Ē��0`C�a����	� [���93/>ŧT�7A@�,,,
�KGt����@Zg�F��ʪ������7ص�9�����[E����OTB���(�U�Mq#�arD|�GYDa�m�VR���i�<?pA����%�.WӸ�#�dR��ٷ2@X�H�y4 �?��EѨ��ǰb�G�n=:���Gu?��<ݕ;?d�2:�J�`����r	�cv�G<�
�#���\1g@���K�����@8Vd����_h��d��~с�GW�ڤ����+���=f��:_X�׍�iB	�]����Ơ�sw�l&�£�j���W]���Y++	�Q�������kb%W"��;��R��fpI%�pGG�bKd���y�IpkE�����R7*�N:� ����G�k�?�	u�beȠJ:�����=���@ⶠ%f��#t����HH�{Odi��A�q�eJp��.N����e�qX[cO� �,r閪]��+�U��o7����'	=4����o��d��B�X{��g���M��db�K
��q��2:��>l���_R�� �
51���x0޶?��?���bώ��:D�~�7r�,�I̳��N�����z
�<fv��N5��6Gј�z_�/L'^�8��kI�\���۹��U���M�oق%E�ԥ�߁��0fe���2���*I��ꫮ٠���N<�`���K"I�ʫ@�X֘J���F^�m;&����F4!f��i̬�]�����j,��uH0��(.	'�j�9V������c��у?-8�XR5�0Dho����gHh�2��?S}�D����X�����!�`���n^�❇^:�c��d����3���-���{vJ�J��{{�ڭ��7^���\~mG.D	Fƽt=m����I�YGv��=g��O����Ȁ��o�]Q��'4�y��4��� g�u\F�S��Ó.CA�w�FJ�{�ۥ5�=�l��o��Y�
��-�B风���	��l�%
:Ac�M��\f�H�#��"�8���c�H�kV;�<�m�(��u�B��4�q�_�D��*@����k�y�|��fT�������׼˼~d�,I����H?�A�ӵ�vm���9��IΓ��jQ�.�A[X����bP�b��u�NZ��:tJTxOH+#�a%�0t5�:�zGs��P��s!5�U�h��M�% q��6�?���^hh���T����#{�bN�ȀbW4�[����G������7�_��G�v�D�����*m�KY�P�,Ҟ���̗�Xxf������"qyV�݁�g/	א S!v+��$ҏ���U��;�-�(�`�X�����E����drRۼ�o��q�~�,�;>�i�4kd{�F�����+I>���8�P�y�%��'��2���0�S��m����!���}���l|H��>�����4�za�kH{�B.��!_eo����`MV"d�����Ӹ�(W0jN�S�=�.��<�;��t�gn���ZC�T��/S;-��œz�+kܥ��̫kO��Bd��u���&��~w���$Yk5,�Ɣ�Ͼwq$U�E��) �������z`�Bw|��uNx[1t���g�M�~�Z�5���{\��%O` m�/����S���.8���Z��S8v�)��L��F��:�!� ��O��ۙ���Ǖ�Ћ��fҼ��h|9�B�:�գB����T2�[}D;T����[�tuE��Q1�V�ٜ&/�b#d��V�{�a;w��o8B�УH��`�i%��;���=��%;'�X�t���[��7^�kᕺ U�����g��	~����l�S�H���V�ˈ���1�9��oۏ�D�;cFZC�,� Ҍ �H��6���^q��������-�����AQ�g��b�� 岙U��ٹj*=W�w#tZM�F� ��3�4�RF	mٷ���[���Vrfu��Eb¾j����epm�y'�09�'��z���Z��<ɚq&��޿�MD���ך�-u�C�zm���
����-t0��AS��ɸ��##�$Cm)*G��x�ZU��L4�C����U�o�����omw<|��/X�TDY������Uub�/ژUV�r�N���'�}��1��R��~QV���Z��&������'�|� .�;�V���F�M~�=K�we)|"SN�#��c���7Kv�Uхhl��g���~<�~�sAx�M߻9ii�7�%L��5:��D�C����%>�n��M�V^���Г�J�	+3kx�-<��W�Q
;,v�)�K\�z�{�_L�������3����f�͇R��b}o�LݺUqt;�X;�*r��W:�R�;�Q,�u�c��V"��1�$Lu�SNdZ���ض���
![Yw@��90\��-�щψ̛#Q�T��ލs$y/��۩�|>J��\��P;gae��JvRL+��X)m��\0�x㘗j��U]^��%�:�Jtδ�8�\�_��GT��vÍ�@}��#% ���Hnx�׋�aD)��4qP�=N촩�|�.Ⴥ;Jh�s���ơ�7��0�Aܯ�"�e�	��s���=1�/Y2�� ہ�����pP��M}M��J�W��(Ækl�x�%.b���Q�=6C]�e��W��5t�t���sD�u�����A����B��j�lqi�g�]��	%"�4���y�>.�|P�0J�nh���Ѩ��.�r �4O=�jd�"�}zl��OI)�h�pGձ�g����|�����{��(�Y�~,�+g�x��@"� m������J�2}E��QB	R�aʄ�	=��=*c�E��6���tQ=�剚�:��C��L�*8�kW�W�-����M�Vr}�¼=5���Z�p��3CN��3RU��GP�k��4T�+&:i�A��$ǔ�Nm����2��n�X�5��C^wu�Y55`6k�F[����D���e/Jg��Y�V�j���~T��!Jzs��D`�+=�W|-W卅x���_Q����8F0]E���&$-"�1$�n���B�_ �v� ���jeuD��Rs�i���y?دz���?wnRn�����g��*�����5�N�8�þK�c����ʓ��'�lPyV�MK��� ��=�{m���W1̐��n\=�݉�-߷������`�D�#�Q������P,H��Pi�1k[�;T�a�0��]������|b�M:Nv�1�¨�ō����I�X�~_;!@H��ή����L�Q%��V���B�y�i�w�^\@��s2���1#�a�c)���`����y����(��	%(%�3#7�@�\l��9�(�V�[�qj2Ӿv��}��~�~�Τ˃��3�@����H�%�U`��k�C��M�5e蝗Xd�S#]� �צ�}WUH̴��mm�$^�5�ާ0`2m����|�E߷�&�R\�D4{2d'9��} ��:��J����Gd����ʋ��FVUL\����h���� 4�u!4�
����F�?������
���۔.f���!�8g}ntFJ�7pJ��ʢ�ύ#ڕ��+4y�a)��I�Ǔ��ڼv8�3ޤ�ҫ��P�К������
��T���}��si�WeG5���u�0�?)��9�D�Q�cq�.���IH�1�'�6�~Kb�Ԣ������]����G�{�+��G�Ͱ�3��
c�q������~{`-���p��ւ�&�9�"��4eyb1 ��lt�C;�/24"c.ols���$��8H����k6�4�t6L���2��J��Z��'�*�M��O���s�Xf��j�2������C�����ʶaK����n9��� ?����w0CK�z/Jxo%���2��m�j�уu���9+��lX8Kt��90�P�n�`�Ғ£U}�y^�\�E>/�U"�H7.hޝ�d���I���E��מ*�<�V.�1^i!�ǎ+dI�_&�Ƙ�\��N��Y2��}�3�����	c�Q��Nݕ�2=�	{�֢s�m�~#ض��$M�����ֶE�j���$'Ȓ
����|���<a�yfI#?��	�P4�Q2�&����mC-�m�3�=#V�5�jh�X���O����?©�*�'��ھ�L�/ޛ��8%��b���:���iY�N��l[�)��5���_�4��[�\�Xz���Bh�S��;]��N��`x��dV�B8b̠q�9�/���xE�=���&|���DD�s��c�,� �� 6�a�c}���a�/[l	���^l�W����:;zU��%�7�Yy�h|�<��[q#�M�J�Tf'��]��a5�l�;��H��pߔ�|g_�'�Ff��C;�\�8'
��$yo�9|W�˙|�$�/停�$��ˬ��>ʃϽK��Z[eL�a �b�N�l��k����_���{�&��y�i�QS��6>':��F�Xt��Բ�aS7��{98.���A�*d@��x�k>c6�A>��J~9�Y����a*��t󚿛`���-�4��aQKu�D{�]*��{Ia�.�m���]�
!$����s&'�I�u.˧��ϳL���6�+[z���_�qO�<0�A�E>��l�>o,q
3˨�mn/�Qxۃ���:~ B�����A�4���W��M>��ڞ��3,x}�j�R
���~9�u��hGi�����5��<K5�x?L��52�)*谕p%��G(:Q�k����#��I���W&������]���0^�C��Bޖ0|]}�l}1��5@�N�����)��6������́��Mn�E;��V7/J(��lV�uv��qҹ��z�1"�[GZ����6m�D��~��o�:�n�O=׻o���٥��|T���V���@�Vk��Zc�:�ĸܻa݊�G��V�Jۜ����I�X�������k"�9�֬�4WB��$�t� Tȷm���_W�<���S�[�Gf*����Zo��#��>;�w�'H���?�+[ŉd����H\P�p��i���/��(9�~@��h����BzC�"~��B0�2b^�zL���K-�S�Lj��4�"ov��a{����Hb��R+�ȟ��a��O�qb�\x�i�x<�hҏJVn�6�l8��6�����U����$���K����Cx�F{��0�dMA٘�'����/l�7�o�L���N�	瓁�^*Y�28�G#6QJ��)�Q�z(~w+$��QB{C'��ߏ��l�@i�42	�iq��F� V[� ���()u���&цHFŤ���M(��^o5�O��9-Z�U�TN�F�Z$ʩm8S� ����w-��UW�ΗU<2�C�d2����+��f]1�	[e_�>�/���R��g�Q�\W�r/,PP'[���t�RU����+��ә��WTT+���;V�n�c��|a�8�~b�Y�ϒ&���ַ���q#��O��"ӟ��?A�%Hv�<|4Sڄ�*m.3G�5�dpO�w9��O��\V�����
 �]��x_�;����#�T�ᇮOl7���i�-89��^܋߀;���~�v���$�j�����F����%�%�G�2�|��=Xx�s0��i��/W�'V�|
(��`Xy��L2�I��yՀ��������f����K�F�	���n4���6�X\���3��~!��+����c�4gE
��%�M�b.�"ҙ�4*ؾ����Ga��-�1ؗ�{P.�3#3>e0t�ZS6�;}�����(�=�D�0`�1	wD��f[ �#Mm��e���4\��@�ӷ?��߀n�[�,�@ ���	Q=\|/���K[���%��u�+����5����+j~@� �S��@'n�ǐ�|}p �M��L
	gn��m�7ӯi��Fk����1�-h��ޏ8>������H�6���ȋT��r�Ki���E����S���x� RF{}L"D0�pO1���y��+��Xw3KmQ���DN���9wt.���F�&���$LoR*��Ӝ��E ҫ�&��m�i���N����N��Yp�Y���s�%x�����Fj�4гIH���:0��NW�\�B�,����kG�EM�F��b*���� �б��tg�< G��J�	�}�;��)�4gg�J�	�;H�b���R8�s��ɰj �/Ib�H=xx�Ê������o�W���ѐ�/�(ذw'�P����:i5#�޼���bY��>�Qq���D|P� �K�.��MR?0�W_�g1�yKm1V�?���2ޘ�u�O#q,�[��ٶ�ra��Ǯ�����ʓ�6���N��[�F�>���w�=���pb�����8�CҔ�z���Ӵ�?��	��p���W(!�f�/iXG�c`ՋG[6N�*���Ͼ<��ډ%�)�K�)
uj�r��"7���@&���P�iܸ����e�ϸS�l��0�����+2e��\P����dh� ��Ŗ����G6�sl�S���p�X�3�9һ��D9��?��0\��]�F���֖�C v�7�?ߕ�m�C�����P�YPպ4���ȇ2�rR�7(��\��Q�Ա��#��&�c��h��x���=���һI�~�s��n=��@U#������.�2�P�Y��)��R��[yP;�K.�/����6׬��
sgs��U��x#��;�L����~�M�`���g�-F�n�"spㆡ����wR�rY,��t���K��`������_�܏e!]G5;��C'�tp'�My̔m��ΎS \4+�+��pC0�CJ�D�a��Y���t[:h[�E��Z;���4׳I��Oq��ⷥ�>�`����0 ��w'0�p�vQ-4	����=�f?�awnl�D��?#��b��2fSv�f�\�c Wb*r˖�5��e���9u�+D�|�km�_e7��`S��3ҳ���� ,���Se̱y7.}��$���%��R�G`�����ț��P�����󢠎���CI��Q�Ak�T���s��b��~�^��p>?h�M\���@� N��J��Ǩ�n\��/%i���W����2U�A�X�W��'�ܷ#��5��5��t�2lMj^��	6[~���UkѴP�;B*��2�Ѹ��gp��W)�e%bX�����Ru�� ;Bf~p��q_�'9���[;�O�)�!����˵�5H��Z_�X��(m�}�<z"��(�T	�U���`e�&��am�a>�j�CNI��?�yE��7F�?a�C�!�{��Dc�W��z�s�%���h�-�_���؆��t����a��l��L��"eu�nHD�~̣����E�m����ۚ+�����q��0.#u�2L��劁L!Abu���y�t���T�a��,�}��Ҟ�l?%���%�=C�Ĕ�\��q����M��ݟG��Zt[*b<�>qpM���h�&U�{���"Rd@��`B�'��� M�ǟ���煰(�E&��GR�-tD�<�m�9��O2k�IG$�7q?�i�G�q�&y��l�K�!��r�=ʎWۤ�?�;�K�O3�PѥI�O~M/�$�U�����CK
4�y��J�ꗞ����r9�������#�R�A��BDc2���r��Z8�$
����|�pR�7��,^C�m�T"%Sdl�B��}�qB"۷��!��û2��ht�̓�b������9�D�;���<Y8�Y4��*��W~���{��)��Q���5m~�"���i�cՅ��l����/��	6C�Z_�50�Z&�z�#�ϑ�8���a%�J6r�*�/O�o
�t�)cY?}b7 )Y/ N�{d����uʿ鄛��	�ڀ��>z�%�m��_C��v����c��N��}�ug6��E�Y��՗�ӫ�y�C|s��B�D\|w�۟�o���fb�9�nf7��4z�~�hr(�,�}l&F������C8�^�N��m�������4t� ���Ro�_�4�ΕZE3q��ė�	U�ybŀ�"������z�C��j��C�+�3i4_\J�! $&t!8R�?U��$��q
���=د��ܲW��:��l呒j3��L#0m�Z��h��ڑ��N�K��<�U�n��w�OR���kEn��9`��c��ڠ|������A�K�O-���i���e�{]Ec=`y�,c��A�mA����֤͗�jE"���jɍ_I�+�U�h�[��)�<�JD��za+sS ��Ӷ�=t��a�ҙ��E����v�7�k"��V�K��K``2�=�{�:��xD��6=}O���smR�C�/�c�~����R��o�Q�����y ��V��]��
G��o����Y�/�w��շ\yL�[�JN���yrH奶�sx ;
<w�\2��J2|��hnAȌ)�K�
=E��xvvT��o���N�`�f3��ӄ�{�-�\��/Q]͞۰�3Κ���NT�<�޺|K�j6��!����t���Y��ms{ι�w����y2(����r��f2�Y��F9AP�'���Lv��T�xom��hġ�,	���7�a=Wʀ`�N��5�C7Å1��R�ڜ��'�Rc  �b�.����t��\��/ԝ��V��"����,�J�0�,�λJ�͐�����I�����s�����ٔu %�hݾ�݄������V��J6��&��|p��^���a@O����(v��x���f0���s	��<m�{x��rI�g�"�*ڠ�W7��h	)�o���hm��m�H�l�U���ޠ"+d�]z���eӕ+d1V�zܥ{X��ٛ7�֛X�*��?�"����I0��WS��1;K��j��u���-�9�cf�(�̌������>�K�bN�Ӏ�/zb�.��שD%�����9�Ƌz�7���y��(+��ӭy��B>�NfK�f�����.��/a�\Rf�JW$ӎ%cU=�T8F��fW~�6@*3|�Cӯ�A�[V�����J�T}��yi��1�+��G���}.>,�Ņt�##���~C{�Sn�l�E�v^{��Xt&|�R��BV��)
V�?�� ����ٴT�oA6�r^Z�*���� @܏�4���������1.\�X�,���ي�@�il�晊�[Q/��gm��n��`�0��� Z���d��ގ�|�|���F�os6���X�f$�eq�*Eq���a��č�=[b�W�I[(U�AS��V�G��ҘUN�In��+O�ݧ�G��wY�JL�V>6���D��Ė\�ɰ�˴�L�l�@9�J	����ͦ�Y�oi���F�una����1fѥ��$YC��Q�.<�~��>o��7Ya��@K�-�]
�}rS�H�4mt���*f$NA������Ph�x��%�)�S?���&2�6���D�og���
\�BUN�**��%����=����(��B��5#����U��_ ��g��7RЭ*��+�R�<�I'��˵6r(����B\�QB/�`e�[�vǚ��zoݽ����1\;�X������F.�Ԉ�dJ�C^>m����vy�G�x��㓢US���1�[��y.l�K�b�gt����z�����GR515����s��㗐�+��D�$��O#P�����\kO�����ￒB� $E- 8�ڛ��?o�@�Q]��;�VG�����?Ƒ�e�t���s�O�7a-��$�C�zl|d��[�㟰�6�D�S˵-��;cx)T	_�����������ٙ�rg�&]��	��z�?̴�U^��� _�L�Ef.���>�=]#�	��:�o���$99@���+mj�>�֛�B����z�U�ذh�2�����\�� N�is�p�w�j��x�;̅��&�*��1������+��Wk9^��{��mBT\�K͵��e<�s���;B�2��$2�'OO{o���t�)�b���w�GE���<�!�'*��E]S�ٽӸ��rCr��8��7���T+�.���Y���i�^����Pؘ+�_�*$�w��n�*��D�������d�q?N�][���(��R��k,"�K-2�{� ��n� ����f��!�߿Ϛ�L;�nŠ�H~��2���1�bUwu�7j��h cY"DpX��1��'v��V`oi����Y��S�C�f��3�N���IÂ�}�d'K���i��I�r��7�~��!^���R���5e���I_h��a���&s���EOzUi1��;���!�q���׽ЎЧQ�X
��+�Z$��D�1��5��TfJ)b&��2A���c�"
��r���a%m^�=RB��o�R���!p�rD����8���Z8H�pI�>!yM yU^?�����km��d�ec��F�N��w�
}H�CWd{�6 �y�j/�+s�+�W�z��$Y� �o9��ѥd�vZz���}E�i��Je�8:&��i�!:���;��B�\���a�=����J�~7%j� PQz�KC��k�z@�� �G��5	��Fz`�3�RԀ�h�:4x)	�����H�3x��
!�.
7C�T�s`�BwR�^��>�>d�l1W��
%���3�`��d��g���PѲ$<����+U��3ڽa��6m�Ag��k�\�|&�o�d�5��O�z'
cvΟlwY�N��{��L#Ĩ��7��[�Hz����C��t�x�ل24j��|KM����0�JW���=��D���Zq����g����>��l��S��0�-+Ip�6Ilw!�^�)͇��+}��w��g>%3$/�E���Ӯ�-CV��+)J`��ަ�l�"R�����A?�]��)7u\�74��j`;m�M�h��/�	洓T���exf�1�T ���|@��{�+d�JDC>��Z���C��n�q���եֹ���Ɏ�i�,4�0�N���Bk��1�HZ�i;Tϛ�~�v?q_�"�PYR(��)�
܀���qJ'A$͔^��@��A�<��`9�'�=�ufGXG�����9���F&7�;�%T��m�N^!�c��ߜ<�'����{[�PR?r�v��O��������5���7�`���ȳ� F��������йd�i��2un_��y�d�|C�!5��\J����m���v��Hʇ���������l�5`6�G�0�y�}a!�b�/bx�5G$�2.��G	��Nف�1�(7���'�D�Vq������E�{@��Nx.��	�8`�����l
�{��ĿG�W�b�!���N�1h�+�Do�z߮���O��s����%��.�#a�2�t&@e9��Yۚ}��Iz/1�+��RW�5|$}���t�@�{+��/�aN���S�b~���T����-�K�%XF�����\:q�E�ǖra�w%�3�Q�"6������\�Y����"�-C�y� ݼ`�N8�U�����M���pCE\QO���"u0���w�d�64�ukv��y�1��ڨқ^�o�ă��҂�#"�k���_�L���h~�O���Q+_jJ�׈@u��AZ}��?�=��J$�dwFU8���%�<A3��@�����h?�i�fk�%Jf�Q�\�G�����_�������[O5����f�[6����0y3��j��'��B�Zp��qgUC�eb������]zl�A��}��E��ZPR��n��i*��g0��2V�D��*�
�S�Ǡ<c�֌1�<TI'+�L���5t�Gy�Ɂܪ���>���E�ժx��큏�&����X^��T���>|�t&���F��Oۣ��s.�u�aƕ%K+�0�:dG��G$Ը�T�q�C��w^��cx�/A^�;���.�W�N�Uo�v�Dk�?�ը�5�tp�#O��*�+�/	n�ϙ�|�*���R�<��%�q�@ճ�PA���~�nfOҢX�?HW���������*8-gv�⠎5�'��_$^ow,>���Ȃ24���a�^]�g��u����j��Y����B�M�{<�Ђ��V��g�;nP� LcRo�z̿���E'�W�~:����:6{��{r�&CS@���"��WR�>0d��.MkS|�3ez���=���A}�V����O��.\�˰G����@�"h��0y�_Ӑ�A�3|GXt�dBJ �_��`4�P��W���à�ply�廸-�� M�1Jl˜^�Z�s=�:����a��qq�#4�,���Uh�P��跏u��(�%�D�v�Y�:x&�Ɵ�S��Z��G�؀<F߽�M�'^y����0Y ���gg��P�3�)138Կ��v�[��Ղ VǴ���"$0L,��d��+ϒ+�H,���~��0�gO1��6�	�-��0n���U��"��8�ΆD����b,�j��Z)����1���=��ݻo\�۪�fn�e�!��Ňrr�s�I���f��	��*�?�T0��P�H��̈́+GjoF������J���,}��HiD�����A�F�?�~P'��GyD�ޟ�F��>E�\��!���3����>�R	a�IwV�Dz"#(?��]	k!��݌�I�����Ba3yi���1�#���Ni�������@�ْ��'���k����^��g&��Mt�ȡ��N6=G��ϙ�45����� ��yIf�P����k�Jҭ�П^�ɋi�L0&ֱ<�D|�1U��Շ�J;�k�88�0N�'���?���,*#��sp���l|ʋ
c6c�0�72�娌��q�5��R��q�b0���.ɒ�m�@���|�l�lw��Y���ΎLo���0���٭.�IAʶ�H���d���OG��0�̟ ��`�dU�t�@��70���N��Ys�n���}����3�|Ǳ�i�o(��&Q�D��Y�Lql�����r8_
Ʃ��>�����v���Mц�e�	$�j�(�ᤃ�xNM^�G�?�8U��ɩ���t/��&/����?�p��������7_�Z��kP]$ӟ&3���"���2�^�?�#�X/x)�*V|���ќ�t9@���k�흗t����@ÚC��_ג �){�$pN�g=E�U�V]�nd�n����^':�<�U�=&��e1������ф�d��V�Z��� ���YUV�.h�����?��,�s>hy��I��\�����$����,��.c.�Mm-AD�J�ޚ,F	@q�0_Y*Hg�
�}�`e�{���,���C'����:gR�|��>�q���\A�o������� _F��T	�AQN{�~�M`㒴�~�{�+�&�q�!�����0�r0�ʣ-�����|�gq��E�"�=ธ�.��tRWH�:ŸC�@�G��E���ܐ��F��p���|���J��P�ۑ���;�`�W�\kě��Q`8���i3�}�Nk>�� �f]�"������O��&>\Y��o{G�K��\�oÄC�ۤ����'w�L}̡w@��k����¨��J~%S��b�)��^�t��犩`��}COKڝ�#�)?4�Dڰ�q~��tR*�!ⳃ�o>j��N��pSO��6��='�?�\s�x��og�*�����^΋ci�E����L������@�{���[����<�B�%�JZ=�c���8f���K���B�Tѓt���8w�|4b;1�����<��8��¯y�G�"���|�{�Ï��xL���Q�I/�FU�-� ��0"�0�2�-�?�~OH���!FgOBΝm᥸�m"AdCvtb/r��v�ڵ���@<o
>u$��\�K��q����s�0�t����D��^p�O�ih5�-l�{g�L��ص3)G�R��ʣ����$��� �Ǿ�p"�����4��tJ
�l祝���}���M��L��^?>�b$�J��#w�Ley+BL�=�M�k�<ࢴ�-=L/ޠ�-�^$��ԥ1��U��t���g��f��կ�����O�8(�Y�7�����)ޓqF!�J���g:�~���&��~ѫC��9���\[��GW��X��%���SӘ����#e�P(���'�0CD� �?�M��ʴ�uP�`��Ҏ�uʷq�y����lncϙZ��N���\>��q>�L�P����n����3�R~����ж���EK�_y�U�)g̙5�q�7����&��ҖX0�����&���g������b�{�����N�ƃ�����=bZ�j>��T
H�@��ْ�܇n:s�1��th�hl!�Ђ���(~Rm�L����}cEB1�����bM�L���I됆��NޖOWي��I���_�����'5�y�6���M��7-���r:�l�{���Ĩ�z�tOlօi�f|�Ѵ���|���_y�����4�T l������%�R6��yT;�7��F@c���
;�J�ȏ�*�D�Q]���j���Gɥۡ�A�	$WW'�;�o�~��E�Ɨ\��R�
z�j�t̷G�����{l�͜�������ά�sB�K�$s�!y�!D����r���[=;d�8��0?�*X)@�_���kE7([$m6"��E�x�1��z� P�b���ʧ
��D�pƝ��A;�	FU�C�p�E�{����q�}b��[Z3��.w�Xdy2�����,ѧQ�Iap�wŠ���_8=.��u��Rf���h����O�l���L��$�Oa��Ǹ��3 3�̌��^S&u�l�	��������6��`sP&�d���T�yqM�f~��K�O��L�eN8o���+�<��/�[5�'z���=�7<gץ{�� �S&��_�k	�^�����[�FL����:zJ7'��vDY&�`H3���
"��_�V�U�)��x>���Jj��$mhnO:Dw�X�M�-���p�)���&l-��*f�ػ�M�jQ�$l��c6Ju;��q/J���;G©c� �g������_���A�����T�NV!m�|�N<���f�b_ɵU�?��On�Xu�]N���\<��3�xQ�x�(��D^L��3Ƕ!�����.5R��l���И.�q�D�a{���0��/�MZ�2�a���ldK`�^L�葝q��ɵ�=�������|R�@�j�HDi�	�*�}�&���Ru�;:�B���16��r�&����' ;�[�J��\5���A������BZV&X��-��
�5����A#;�II��<�i���=[YN)���ѕB2��1@�>�z��u<�D̂�Y¥;D$U B�6%���p��)u�d��C12��,�:G��lBܽ!�f��u�/w��ɷ���Q��+=���j~T���M�7�W�L�]�~H� -O��J?|@昢�>�]�L��PjI�;-)xZl��T� F^)
1iY)���y���%E*US�u��qd)�Z�S����)�A����H����4�E�/Uh7\��8ur�u��p4��;>|���@���F Y��[�\�D7��,C������9�8-\�L�b'�4on&�ɵ]�O���7C�o�{T��³T�U'�'-�ᆶ��m[:����Y��z�8��36�#ф�r�Fܵ�n��
rjR����Κ��F�/��n���[�Nb�o��_�*���vK(��m:��b��������-�
-����\�o���0��_a�3�7�w�^��3bП��~h��x��,\�?� ��@r���P���Em�tǧ�]�uØy��oN���l����@���9�1�}������D�
)ׅ{�d���2
	b#���yR��cf-q���Wz�k�xx�Ȱm3|��X��s�b��?J��TR��@���������=�� F?��r�eo[l3�J���P�z��ejR��bY�¿*OD��g���E�qIh��Sɶ�z1ȀU�>~�hH$kXu�4^��F6	@B�녊e�%�{<�g���e;��Dx�!�����M�����Zo#�/�g�f�z;�g�L:�פ)�;�C��gq:8�e5;i7���4=7��:��sO�s���&�޳�!�Ta�i�p�}Y�ha}��9����uA O�p�"c en�>����*�W�����	��:�%����MX�Rb���\1�-'�bSyX&���S�d�U��Ƀy�R������1�@B@$�wq�f;>�m�5��Dߝ������UO��0r#����b�r���f�8�̑9���yZQ��~n�2cc�y ���8�H��D-�߈���JWu�ý��&��d��w	t�%9�>4�9���yݽJy�ְ8�s���F�A����h%R�O*t7Tv��I�X�V�;�gauJ��,�V��hw�a�v6���&t6�4xPע��r�Vl�<��t�^ l&�"5v?x_��l��\�+�S�k��_���5�.�߬R!�-ңMnL���QͩUP��VY�raT^ٯ��3�D��&Ԝ�++��Ğ3�&��q�"�k��4�ř�����$%���Tl�RjW=j���a��^L��|RA�xY�dy�L��_��u�oX4���I0��Gj�U��#�C�.u����zĞ�!�̘����Rw䞂�k;�J���|_L1Xu;`t����������ȹ�x�vTLF ��4+I���ʢ�������8���f��M�"b.cj�j��*�0���#1�������M��42VCRC�h<ܟ����W˽*;3�g��'�h '}�=ߦ<�=�&���j��^�I� W?�FDA��;�JA�6����a?�3n9
������L��Ũޒs��wELa��Cם�]3V�Ϋ�%�_�g{S8`Z�xQ^/c�;{.,�}�m;�dj����V�	?Fq��l���機����8R��Bs�Nwq{��o����
�4��S�E�"��>?���p�Z��x
��~g~��i�f��0Z��P̠Ȅ�qNf�"C���X�����$�D�^϶&�iN���� xȸ�h�p����ě�9 ��Zfe߭�?�� z;?.i+�b|���+�>Wz2���4`X�'a��M�v}ŜG�c��Rr)���'B^k��`'o��-5��Ǎo�<�z�gyq�C����9Dx�4�H�ax���u���Ɉ?D����?Qs��/0��&(�Zk(����v-��8#ɳv,�ɦmhN��0�I�B�w����C�rEfo��&ɭ.������IdB�rRG$��\�T�������J�*`S�������j��QuD��A>Լ�ئQ	5 5F2���`~�k��J�@�c��,�r~K��
�ww�x�Aj`R?ąb��%������QϘ8Ik��
�@{d�[���2t�p��Ʉ,��/�9��l��i\���ښÐ҇�2Ts0l<��^w̳��[����pΤ� -arr���Z��k-�^0�Wu����yT�� X���_���I�E?`���<:��9��§	����7��զ���
О�����x`�I<���@����:˷n/̠*��rY
|�D
ɬ�����8�O��X��'��A�lZ^�fy�jD�H6�cZ$2>�>,�Im��;bK��UwZW�(�|G����?��l���A��W�;��z�m��������Kn�/k���۾I�t��zV��jrg�%sp��	�}&!ٝ�;%�1�[,]�RQw�>���o�wnļp��ß��*5�K^�o�|3
���W�Y6��x�x��ό�~F��j����(�&�˯u��j�%!���PNr��*�K�e��r�gY]/��k�aXq�r�s��v����ş��"0#����ף��]��ڇ�uGky==�^�M��؋�� Sû{{]�Q���%�k" ��}�M���w� w��&Ͷ:��>���hщ������,���K��l��i�K;e�=�D9z 8>�c��I��𷮴�%�m�(<���L#���q���"���C%f�����KXo`�]
)��Y^>d�C�+�����4�{嗕OVS।��j;���m�hN���
��E_C"{��ϝ��U��$�^O �8���35 6�.�a�8H�%X�=Ȋ�MgU���x�v�#�����b�	!P�� `*� �4����*'�����s�(�R]a��W+x���{�YB����R��cS7�¼oґ�Q����Us���.4�$/[t򃱑Z�j|��ܤ����Fh�_��ا~�u*������UUY���Ģ\Mฮ}��7�BM���}q.�<B�? ����KL���];v��-����'N�`K���0�\g���J�eM�6���Df9��7��)��S�[!� Ks��m^�����b�,��Xw���'���/���0�ɝ�{�'��*c`����~�O%S�9��;�q�Ӣv��tno��}z����y����ИQPK)v��P���SHm
����5��Uܺ	y������?!VI�϶�0߉�lt���9[�T�qƶh.��2���`h�0klhM�k�J��j?��d���H�J,I:�9l���_�z?���1�r���Nc<p�ni	�[�	�ݛ�*+�4� V�ǲ��B�.r�$�
L~(�~��l↎(�:���&Q[��
�(����k��멊dZ�J+�tF�?��֞c� �g?'}7�a��0>�=���۳�P��%ۍMv ��c�m޸ɥ��p /E���B���˺Hㆺ�:w*���l]MʜS�_�@��0Y�sV��(!����Iw��y�e(|��6���t�����J�q!�D`��;��΀�G�]�7�N�3KM�@���3�R�}H(��(σ���ӗG|W�
J2��m�߮����l�N'�ƪ'��'�XZ��T���t��٭�x�~7�;�p�$ u��Brq�&tOŷ�����l?a���ߖ�rƃ��!�˗L������x(@�?�0����/��T�k�y����n��򚨕G��j���6����R�'9<w=:�<P(�6�.��~Jb5��FÙ_����L��>��'$�P�4�q�_Fī�̅>�A#B�����{��߸�l�j���3�WQ�����)�lec����;!�8��-&��J,z:)�C�U/��7t�Kٷ=�&N+��y��~�'�+#>�;!?
�7��h��`���A�;8�ˀ0���'5���?�I΋;gx/?��, �����Je�TF'��,�j
`����Y$jD�ʉKOZ �CG +�QcE1����kb��Pφ+3`�x'H�p6�n't�����铲��c)pZ3K|�����SG=_���S�+pyѕ��ɠ��ً[����epO��>"վr2�� �,;��������,���M��-TQW[�ǟ�f�0`��a��5��B��,{�U�(/K�1�����\�
�Å�����4>pط��3��7��?��c����\o#$�9�6[x���M�tg�&�G�H���"�ѝ��}ϤG�*Y�*b�M���~�2�=zyЫ�!�	�1�B��:�������Ԭ@��Y��t�����^�UW��f�#�֛�y@7��+d����]���	$$sf�E�3�0e8d���Z����<ׯ�Jz�(���)u~D�O擓jC,�]����4���j=MzZQ����ΕJd��:u��<���A�!G{��t�5��1&kMAU�O��������ϧWZ֕`�8EB�Co������[J����i����r� A�!3�Im%��DT�|��z����J��(�Ȝ(^T���Jن/�sI)/K��� * �f�B� ��C*���ykZ�&*��"�X�YS��o�+V��rpgE��*Oͨ�g��_�D5 ���~�����o�o/̇����ৣ8,o�ضh�Y�!l;o9gq ]�rƭJl������}�m����<�vq )�����L��]7n,%=2�?b��ƞ{Ʃ񎵒��!��@����� ]��1e��TK���Vm�,[4���.8������ '+&�G*��.)�5��nO3:w!�8(0�$��II�6�zkc��4K�@�^>!��lP�u�dY��	q���
�+�{�	� �d^U��mG�u�o�^��$�Bej�v}9�e'���902��w~��I�2�s��#+tF��������|�X��8h��ީ���y���:��7ŏ���D���{��u��k�H:����=��AU�lr)>$�>b�8��Ɓq����)���O�ޏDl��,լ*�Lq�j|�g�Hʹ=�c�Ǣ.�s�h�����x���n'o��R�Ϳ��on蘃�4\�#۪v�!�DL�r�O�׼2T ��W��5:�+���ngt���R�T��UB�Ө��2�J���`��mŬ�� �XuU�~Խ�Ԁ��L�r��D�[�`S�d��I��2rk!� ���ϡz⿰��%�6.M�E�rq}W*����:}�w�C]�n� :Ǹ�Jd��������8w�Y� �Am9'�!��\������g��_̲��{8r,z&1���Rjc�n�yq�����F����>���������bNFOb��fvkB?srz�| �.O���T#�v4U��ڪ}䙾}H6St~Dx�9��[v�^�.ć�_��fWQ��E����訰M�'��,ͦI���'	��yh�����v��\h������*l̝�q�����{�<���Vvq�P8_}��x��>��e6�o�׼�|'���ѿ�� H;SLzSӯA���s{h�t�iGի?����UN5P��x����N4�Q���d�M�
��iJ�-���ti�Ț;�G�q@����B�aLr�c��']���Z��@�ZtNb�m Z�|�ғTc��|���ǳk�6�7u_��a�����j����3f�=��b�/�h
f�?��;��#�JK�;H�M�[����d�/y���6��M�3i��5�pY�o@c�[���
S;�K� �o�D��?}�WT#'�y���i�j��&�����-޻O4���d�g���G�^��
�"0����#���
ŭZ��|���.�)�$&LbT�uP��;���O��i��󼷉� ����4x�@�$6��M�&�A�,(XcP�R�����P��|_����K����P���.��&V�j�l��Ȯ�K���&l|Jr�Ѱ)��Jfe�ю��I׵����iГc/��y��-հF���<k���F����@�!U�x�~ �B�X���>Þpd%�ĄVQGp����9�v���G1�A��I��e�vC�Ȱ"4*��B�L��z��[���Ё��9�4 U��nD'�w�HϬ@�t|�f�OD�v1�o	�^�b�(�v��������([
Iݱ��>�\��.:΍���W��:n-����grW{d��Mh�I�MnP9�G�4����RA�Swqo ���N�uj��c�}<��h���*�[��|�Z��%߁zg7���z�ic}v�~�r�(F��F�eѥ�?�M�F�V]@_\^�gU��Yu-��}+�Z�Er؁�ڛĩ8O�L�Z��OY�K��L i�Nj���S{GYH��h�ۇ��]b=�T �l��JGI����A"�oщ���t�ٮ�� �����+p��u��?�^+��(V�+�N l�О/:�`w:��X덷��08jp������P���cq���"8Z��X$���F�Z�ǰsx��GX	2�"���"4��L�]`?1e���S(��o��p��jp����u�4�óHm�Y�oƎ�m�>�-��W���y�h��s4Qt\"a
i2��a_�Q^4;���jg]^Vsё��_��Szx^��Y0�{ຽ���[R;JW�C�慯Ҵ0�\{Q'�u^��up�<0���}�[���6�,�^�1Ij�&3C�" ��"w�=c���h]&7������ο\y��J��|�K�#Կ�;��]b7��P�r�\	/�1������<+�+W�@hS�bq##?|�����=yf���HLpZ�qf"�*8��ɉ����0���t����p2�F�
��0���/�W[��˜��(�'BG�'���F���!}d��!5��D:��SjXQ
���$��g����4�t9��y�"+�+@(���D%�12�Oޢ�8�Pb��cP���t�Y�J�e����Vx����[B��m3���IX5(Y���2���9�5mj���U?��zKCXz���R{;�3���Kq������2���tqƱ2�%w�~����SS!��!�ťtz����,(��xQ��`F�n��jg'1��3��2_���Cތ��\�=~��. t��P�Z�!;�?N�7Wܪk�7%W���Uxl���-0�Y��}�{�-\��]��:*��j�d8S*�Y�x�S 	�	�pj�i�<�|�*�S��U��3�SF��U����]{ӗ��/X��ű^��^��>�dސcx�$���Jষ�YG.�?�i�m���8��
���B"�Ҿ����������&����[#�b�o`��uЇ�{;WPǔby͠�F1,��m��竾�+�8�6Pc#Z���R�|�r%ሔ��:U�l��+�fhg�Sr�SZ�� 1�mj�?p����yڼ�\A#�)��Ge�C�E Pb�������샆i�/T��
���ٯ�r�����hs���]��):|����U����Q�o*����NO�ly����T�5�6�^�lٻsƺ�󇅜���,�Z�� s��g�;b��ʶ��i��NW�|b��*��d�����M�VH3����s������22�,��P����E;��}��8�p���$��u��ၕ35��c������l����"���޻; yWi��M�}�ɼc~-�/����ʃ�#)F2 �IO�!N"R�ݮ��ɸd^<��{��r�H%L[�^F�!2�y?o��5��z�&�o�Ԣi��P�!\�k�.��̕զ��B9��i�w��C��(dz��p
&��X��`�g�H)j��9�`$��~�iׯB6c>��~�/���QPa��A`E��`��&��>C�25oA��o�[j� p��Ԙ� �/�E ��+*���_�X�iI/*�NgƼ	O`�ݐ�뛏�}�W��#�C�p��=����0�f)��U��SQ,�I閥!�EH%=r]�Ѳ���D��:d�q�#D���� �" ~�)�`�([z�;���B-�Y�L�7��͈Է�7\kYb{�4ގiٔ��@h�1�̋T�Uq��k\�j�,3���[V�Bg�2�V��Y���M��������^c���!sK�{U$�ϙ�rk2�Z�'zm���3~a�����?�|ȗB�J�%�+�w~Eoޮ�&���d�*��D��=�%?e�$U��|��'��+s�9{��$��D@���"�0�R]�Z����sϞc,Wq,�}ع��{I=\`����%zJ�l�	k�>vԖ����<��YqW��)f���ZaOp��D��P[N�	�Q:,���5����4|dd�A���Z
j"LҐu�m�_���Aw>hrl9��Y�6�[�� ik���p�"��q.'��Zrv�k�5������&��yź;��v��-����E����Ga��j�;�VM�+�#���7���Ю��J)�}�� ���s�{��>vP2"8��{ֳ���!5����WpA���ъ+"q�ޥ�'��$���*�9��@(3��J����֘�x�"$N����<.�nN>?F%}�Up�gU���#	��ð��X��P�'�p������5 t�&�$Q�7����"�3�K�^r�辻Pn�)^!��U' �.U��3���_dv痀�OX�T\lX�4�5D�3o����I̯�/Ĳ.N�	s_b55��xj��e�hK��7Z�E������[���C�.��O�Q�wڞ`u�=����@�aN`�� �Y�Ou�$��~��ױ�u$�3�ᾎo�v���HV6�����p}%8�T���K��Y��=Q�!z
fޣ�p.d�9��wm�4��rU������1x�xG4_��;���`��YJ�T%�����䗆:�08q�Z�����3�NYKz�!��2;^pbS���<�Xdc�v6=H�>!���.�7j�T�����J�9.�*{�%׭���p�����j6zyW.��yW'��ҥ�2� ���z�Pߧ��8|�\���pȜh�E�J<BDD����u��1�w0�ˉ�/��b�d��PD��y�-��ݜL����/J[=�F��Qk��Q�8���.��7�r<g�X�4bz%|�7^x�������fuș(FG1�����x�@ό}N+���� ��@4�8h7�Lh�l�v��9��5)����#B�;��r<�,Py�`��z�ĩ�/?m���]"��X�6ZzVϫӓ;��(�=��]2�p� �"N���c�Z3n�>(��jٙ�,^.�Ϝ�{J_����P��qs�����u��Ry�㳋a1��b��&�ݚ�l�	=[���G�i� ����gQV��Uѝ>P�t:�=Sh��4<�c>�w/�D�!�$��P5����lp�G��ɶ��ar-�`�9���3V��UL`ZWp�'�è��X�oD��b�U���N���_赏RO_��Tj#h�/ɧ�����h4�-`�X���[K���}��ehA���%��c����04��RG�@���s�U��,\�5 � ���zoΎ;<��y��jZ�=���g�ֲ�8�܏�@n�ʨ�MR�w��:%��|�>u|"KF�i���}���X-�� M�ŀ�A*I�@nQGl��1���D%������b�������G�J�#�Ǐ4���R#��(I1�i����r�F��N�ZԂ�|+���0m=-C16Y
�fꁮ�žW\�$,�X�P=��y��d�����Rq� F����ѓN^vvA��{׊cc-����I]ST�٧�%'�ć�7	�W�3����R��r�$vZ�����	�-"�wQ�D��ž��X��?_0G��*�ɑ�N�l"O^�A*3�H�S:q��M0�G��mK^���P�\�|��ئi��� ��W�"�wK?��\WUX"�<o��"|@bx�Ж�`cD��^
/(ñ��l�E�,Ν&c<}|��������)qƴ�MA��`����*���bޯ�����b7��1�y�2,
�D�6L����}�K����r���J6z����Mޤ� ��\�y���s�8Jt���AҘ>�ĩ\�Wp�8ǚ;#��Ըø �����i� /�G\R]i��a�`<�߯��۷�	D`z�!�bb�f��E�1��%[B}��=4ܬu	ך-�*���4C�w#��.?c�۪Y��F�4U��ժ	�U���z�6pN4B�MD簝�Y��5@$�fw�e������l;�ϯi�sQ��/��ͮ�/:n������[�,��	EU����A4��[�J���˳E�|ۑˆ��f��ꩁ������4{��0�ڏ�����$.��\	R�k�(�@���r��j�o���XM���9OMݏ	�����%͟�4�|6 Ş�#綻��FB+U �c�	R={����'@[a�92
p�K��Ψ^8E�K'S�����s�I��{uB��2N���M�dmEt&�;w#^'7�'�(�h80Me,11���NYu�'�5��Fum7�&�怙���OE_�hsK��}P�>�P�V@#9N)�Lu?��cjK��ωA�RW��ۃJ��R8��p�T�2���	46����ƃ��l�
����bX��ֶ2�gH]T�
����?��w����r|r;m5��ؖ2壡�g�lX���;fc<c�jP�t8㾫��+Y}S��r��+�uS8H��7��[:p�1�+��Z��t#�!�����^��I'nL��p���B��Nj��fM���H�gP `�ߡB�Ueu���)� ˰�\O�~�����t?	�>
gr|�o��?ė=�I���\<�Scyg$p� ��(��.���tb�q�7�UKZ�n�RW�n�ͧV�����	�ݡE��Pm����~��C]�Ϛ�G��0Tp���Īr�6Bh���P���S��=��dA��
�·��*98���z�v(��>.`>ұW�ieC��e��gv���=�W���ל�] 2�XWw\~�}��&�����x9e���o��b�ݖ��s ���3�䳈���%V���fQ�K��4�JH����6��S_.$	�,4Y/ʙ��<~O�3�B�w�����ʿ#?�;̉Pa[8��B]q]���7���pJ�a�Q�f��\����X�#p�c��p&�5�k���O�����K�,��Z��� R#�0��o{>�W
g��
�*.JqE��G��-���^�q�3�v�ȩP��
�c�ꋋ�v���.qӣT@��(���@�	��J�Y��:�3�u(e������5n~���̆+�ҮbRX{ޒ*�5Ix@� كT2_^f�Q~�t%QaqF�"y�˓���ѩ䙫.#��"}�oE8P���Y�F0x���8�d�Ɓ��kI��p�Mٜ�W]����fZX�'o)�#�!Ԙ��o�4���\	��5*O�L�FE#��
v/fA��5g#>U9�[�y�{��Oe�a��U�Y�@?,@�(�$�{�xx/����9w:H=��ퟞНV��?��$3H��W��`��N6 ��K�f��|S��[��ڨ.�%��f���+�0�_�Co��S�F##��_�fL�3 �V'=��:�|����Do��ˮ�#���Bgl�U�����y��3�!�?䏆s�ٳ��2��Ǫ&���r���}��He�eς��N�~gBLj��$�N>|`��$�V{�J�P��w�Bm5.�1)?k�g�&i�v�_�����+�<����o�Bp�*�0�s"��	{�5�qbAtK[��(9>W��[���h��̪L���V�s����GW�W�1i�b����)ۅ�Q�Flˍ\67�L��F3�[��^��x�u���(B��EP��L�
�`2]g��F�T|�����U��UqRЅ�Ҙk�mY��^zU!�P�!�Y���'(oi*�0�8�R��v�ꆤ�r�>�Z���FG�l���"��ҧ�l�k���1�L��0A翁U�k����j1S)g��T��؊ ����U֠cA��d�+�ȀF؉l�+� v� '%�ԗ�-��㯩T�O�3��N�"т�}�å~.��r�r�dY,I���u���VxU�0��7�野cL��aA�q\��"��t�)ݦ]�cki ��Q���#Z���׵m�X�_�4�ø4F0�0���]T;�fc8�cx_@�g�fu� �y~���$�͖�/m"=a��E ���u�):$�(�M���m���ۅ�����~64d�������H3��;�u�#����&�P4 ��P�J���R� A�2R��o�tկ�6s-:�p�@�.�ۓD�`)хc�ޤ�ւz�	l��0���� �2�}��������h{�5�<|c�xs���J�Rt
	��&Ph�>�Ao�#l&��^���-��w|?KƮ����_�DKq)
���0��b������Ȕ0�p�H�7�~x�XQ8�X���f#X0W�%�l��:q.��/Bc�����q��-u��,�f&)�bZ|1����sdh)m��n-�c�ex�P�������]�T���̅��]$?��>�2?X�ʗ�~k�ޘ�$g�Z����LȂ;4�x��M�2�t��Ң����Ov����΅ C��[x��,d2�s+�U��d�8g�	*䚨4�qI��p_�A	z�d��Z?r�[���=�} ���܆����C��K�H�P��C	y$��85�1�~�7�i5G�ݥ���>�Z�Z��A~H�7w1��l"r3�ph����;�Ҙ��6�H?����� �_�p2�y`)lr<�"�d�f׵	���K,�+�N�ط���:�I=Ӿn4q{o��4��+ٜ��:��{bӁ��j��Q�9����UZN����Cɾ��I���|��18�W�WJc�Ń-Ä6����r��!��os�wd+Q#<^���J�]ZA8������LExt�O:���H
ڂw���k8`~�P¨����]
t!�M4O���2	i�oR0�o�����3�L9L���/�J����b:�&V�z�(7w�i!]���~6`ԍ����7��2�5��AeK{F���I��i�)?����a�S�Ȓ8���-��BF���2w��&���d�R۔���	���C�t��)ƭv�(xB8� ��$$ۓ?���Rb �u���Č��z��uM��
�%@"�B@�a1b�������\*�~i�=���S�I����ry�wf-�O-�'� B���v_�1�����t�~�����K���x���s�j�]��`���l�����3Cf�qbuD�b�KG��+MML\]�Pig˩4^U��f�E��.$jl��v[ғc�#�F�Y��f���9�1�E�5�ޔ��֬$��<�v�H9�eb/�>�W��<�;�P�-f[��t��N?:Dϭ$��s2�]��A��a�hG�lD��qk�[:�in��Ż�8��vj�/R���K!��������ퟷ�R��ĩ,���v]�s��;\6��m$���� -��ydq�j��/-�N���R�6'7I�����Ч1�4I}�o?c8�<���fx��rm��D}#6����B;gV�M�C�!�)�2��7F�OjNS]g��� �W��ѩ�hڈqԘ��ѩ��p����3�)|��[��1�AqN>��Ԙ�A��V5g�I�_� �6�tQ���[~���C��#̮߀Գ����u�V+�Gd��j�a�T@}�|������,�OA2<3@�nc���=Z�j2�Yq~��Q�sFxP2��	|��B:b��D�=�����6�>�!0�.�����c�c�㨫a�Ei?-�נ�GI��|�l��q�Ë.&6	E��P�SP��'��>*�� �A(��K���7�v5�G�����:4��/����#�?��lHx�@c�<!Dz��U����3Շ/J���^�2��Y��?� ?(�|���ŷeD9~k c�Yz�m��k�u��r��״7?��.�I��mz��wk�M|6��8R(�0���E�B;4����2�f��G�;b� +�T�^
\��8%�� ,"�xd�<|#�ciN��)�-��(��_A��Ť�l��D���穀��$�r���pL%�Y]uɫ����dl{�* �\�t;�����JV���[�z傀n�7��v=�'�YH���o3��u�\m�kk�CΥ��
t�X��-!���M�ۯ�"P|��E!�b������� l0"��,9�D7�W�?�|*$��H�~���3�*��a�"`��D�&�*B��ɕ��.Rx�2:������e�	���l�K�$�O!`%��qqr����ٸs���$�7atiG��4�ؾu�d1��Pc�z�	�KWbD�y���M1q+K��y��O��˦��U�ճ�%��*�P`㿅�ь��ɰԐq+jl��ChR���#>q�J�L.�%�\/3��g)��V�5ݷP=�.Ԧ��mh�!�S�Β�߇B2�1"r�
?:8�9�܏@wQ
wTRzl޳�!6�Į��Ȑ��%�?�:��S�3j�"��xN�L����:�"��^��Yq��}0O��4j���[Ǖ"������Z[Jw틞7z���z��Y�9:ȔT��ޝ���w��R�=DKJT�g�����[�t���Ѫ��4�Ϋ|9-�_)��1��8
&Z#Eok���<h�
f4�ᱵg���uA�q�DF�qz*�9�,�a���%;=2e��`>�D�cOF���Y�ͧ#f�"Kʣ��_A����7�@��1ť"���s75��E�1�l�<P1T~�'����
�|����2��v]I�#��6ʦp`,❏�}�	���Ԭ9W��'��
��n-�L����z$����W�t��Ě��	����ÈEg�Pj����s�*���S�?*k\II���u���dOS@�b�?\ffQ����)�F���/���08�I_?(�q�Շo�&��4��5o�1���W�������]�A�$�rX�lbCUk������V��ȡb~�HyAkڀ�r��@$��8(SG�1r�	.���xF��Tca�R���t��&'i�IY�08��s��$�/SJWP����E(�{�ɘ'��<"'��4vG0A�_��Q_����+���K\ʘ8���� i�ӟ�B-ճ�_�r�0��B9՟�Ӎ9�v�������Db��* G���tEŞBD��T�kY�L�H�h�F}]�i�����O���+ର���mf��UA�;���:�v̯����8�x��4f��{�2�K`O�9��Mp��B4�1��iL!�A#���OE�4��Ġ_���v ><q��O����9_Y���ioa�9k�M���%�-z3�幝E�:6�r��(蕧;o�!_��m����pu�^K�b��4#~,`��ds�{L�-S~�N�`!��:g{��,����:Ye�/}���&)c��w��{
h3����W��Z��:��U�O���,f��PU`;�N�x��fJ�~ʮ�b�0ڐ��u�+���]�B�:��o��?+�-���H�hX#������j�s7������`
VX8��5a�񬘡�:�����谆�Z���UuNtp���Nۚ��bz%�^ݷ�}������(R���$}8}Л4��t��d��%vN���*���%��*,L��S�� �������l�7�5u6�im��Z0������{k{j�m��K���<�����:�v^FO����1$����蝝���@���]2"8�⿯��QV�.
���U�eQ.w�ҙ�dU�|5��⏌�~�/Pr����4����15���=�w�F��ɪ��1�z��g���PH��}��x����u$�&�ݪ<��g������Чg�,��<Qº6���I�� �M��4�{������h�|t1�Ô*���7�8�M�Y�U�j�		��Ͷ���*L��a��5���~ ���O����bK�3V��s��t�\祭��)08�}�f�@<	�1�<@��%�N�p/�A�c?&p��ӵj�Wܘ����eǅ�z�9 ��Nٛ@��J�ȅMԇjD���PB��^L�i2.���,���g��~��$JE=c�W���_��QӔ�%=n^���ј��9$��q�d
z�`�Q.g�F��;�H_������A��Ϝݙ��.K?����$�' q[�I�Esf�1�Fb٭$#s6� -y�1�J��G��#bD+X���iS���w�?��>��V/���L�d ���#A�Lo��4_�I���L8W�u�lI�/�x��f��'zԼ�HoP=7�9�>�ѥ��>�Q���V^1�]f�,��5=H�z��~xp���lÿύh�~㩵�s!f���Q"o�H�8�����hY�qd��z�)z}C��(w!n8q�H��*,���e��2{�Dz�&�F:���j1�濾1;��L�Rs8dmtQ�F��Àk�����},������sc 0J���'��&Ga4"��6O�XN�=�UB/~�y_�M�S{�7�9>)�����J� N�=m���e*�w��`�+|7Y�JDz�G�Bm/�sa����GSX��P���
~=$�Z��S�GA�x\�,Q�طOn��:�<r\���H3#����@�Q�y�A��Ծ�WF�SYD�c�h�A�CǕȡ�m�����TJ� ��([�&�!BE�� )����МJ(�Q��`�TqR�d!f�a�F���/׉9���-��e̙l �|3�;��I;�Cf!?�{unAG&��=2R�<j��!c�%-�Y����w/�xa�u�[��O�)?}�݅�����#�]�eX��G9�Y;�^��|ٻ0AQxm��Ը�	��7��ry�!;����
8<���oV,A�I�"BtV�R��Y1���Y�������rp&��W�_�n�+�O{�������Γ
�#W)Cl�}��LƯ��f��C����}{K��ޙ?d}<HM�R�~=e�D�L��J�� Th5��g�nǹ^�oAI*��-7ᨿ\�b�Ђg9U�adyl����H��kdn������d'.Ǚ���a¡��(%N6�EXN8���b��x�h�Ki�Y�Dn:���,�&f�0��v��zGIa�O��H_C"�ZI��M�Vf3ϡ���aT���5�4Q\Dނ��F9y��=���1��$�B<R�PUS����+��0iX�+`5p�����[�����ś2��Cӽe{�4��	%��5�����څ������|-��^��񁁄�pi�-0�gTW���^�D�����M
��h(:��0+ ������?]��IXO.4����!`���w���C��ن1�:O�Q��Қ��yk�.��S��(>�H<z9��ṷ���7�@�<L����4��C��.\(����\�ʔ �>/Hw��I�c�Zc\�o�xG�]X׋�4��c�ஞz�o���B��Og뵂�)���������R��� �꧛ƕt��Z����3�ZD'���]�祀�uh��@E.���zl�HBc�A3_i�z����[���!鮁�b��mS�K�N'�dv-��p��m�9�/!u3�dP7+��'ƂS�S�Xv 4��R�"=����R�R�s��~����t�����
�l�n�έ`둯������F0Ⱥ�z�{>�f�bZ:s�����8ѳt���륟�^�
�1��R���s��n�E=��譓����ś�b׾��Y�x	�$���E�,U�W�"e��Lf(Tv=�7�R\��7G�A�9�VLU!��O(P�����FU��K��%�/�l>~G��8�X�
�p �T�aڳ���V��w@�VA�<�w�����9o�5�	N��>4� L���:��貌j�?��R^���]�ccV�IWw7�5�c��1?o���:��a@�����#�?�)�@��>���
a:���;f}S4�:e��N�Y1����0�~: &E�<M�����s�V��J�2BQ������U��wH�i�H.~������ė���ف����Tm��A*6yN���>�)=C-X(�����d.��]=� w��%?9�]Lvn��y[��#��c�J�ʉ�4ʠ+��f
f��V�O�ykV�
�C�]��!�I���.i��^��U<+�&!�Ȧ��@�k�~�����4R��^��-��Od���\�za�̫8�J6^!�j�oP6��&Y:c)c�n1�7,�D��%�et׋�,��s����������R��M��*���ڑ��.I����3�����ߧ�|���RVW:�"�q=q]�#'�+��cs��S�UV�Ǹ�Yrd��aj<��Cyɀ�Y�U�io�4��'؄k-�Z��]h�^��`t�"�\��P���|ơ�T@a��U���6}��ä6ڏ�E}'/7 p+�=�Ag�E�H'@\�l���!qO(떀]���L:��B3�Ŷ�%����D�T�Q���F�"Ku��h|��^�u�6�0��lcN)�=�i$�ݹ;S�?/Eb�}+�w�?m ?�� �^������3�̽*��*�`eT��F�����P]��
�Wq;8K�%�ɕ�Z�nJɩ��zu ?g,���Y�KԎ\|q�F� .�Ti1��D�G��\� �W��e�ƀ5x�k�J�(��7��ó��+��;���To��k7̌P����x���p��}�=s'C��R`�ʎ��]\d��oE��v�ۑr{���Du��TBI������yX�[��I9���F�E�]�vۑf<�\}@���_�*3����I��|��-���8�Z������q���;�Si�2jR�����վO�'�*���I J�(*GX(ҭ�c�O�#��_h� �խ���勵M��|��3ݑ����r���
X�adY���O|�ϑ���" B�����Ŷ�_�t�W���e=��<ε?9Q����)�$�T�8�<�aip6?0��`=����}A�g��Ox�.L:ƍ�>1��rH3�]��)F���Dr��@Q�]�b*e�|�"�g������כg�� �q��T/`��6F���/��]~�=փ��?'H��]�r$���'�.+T���hsYpY��.�!=�!5��5W�7���9j��iY��m�ځ� G��Zs��b�ьLQ�1428�
8���M���v��O3�ؿ��h����L��M�'pA�&�P���P3�0�����F�J��Ų����B.p��CM���16'�8o��!��ɘU� b�'K,���[R��t��rPR��{���^��ގHw�縯�a�-ۮ"�$'O�f��@(C(T���uݿ�@��;�P��/CHc���v��	I�ӹD�Mg0�9�W�$$��6�x�y�
�n�?ب���I��έm�4��x���To��U��o�Ǯ��U؂��)�dF�������%�\|`�O�`����<� �4��yO�����rq����r��s����G���R�@��-(`�K=��T�2�.[u�+)��4U�`Q�������	`�:ʫ���@��z���W_�%�O/�߻=��#��@��q�VB�0H^sD������YJ��c���n9:݋��ۡAA_�ju� ܺ��S���9ͽ�	�\(&dZ� �,�w�����H<sI�m��չ���9B�}��[�<��&�.��Ӱ��  r(�[C�����ӹ�1XW��m�I�.�|h�+Z��=b� R��??�f
�iF ok�3mC��$h��)6q�3&�%R����x"�{E35Bec��{n����B�h.5Z�C7N�M�a�=�"W��:�>�ɹ\9��]ʣ�n
�����l�G�Ð��o��	V:��o�
d��Wld|2�k<"]e�Tja]�v�O���!`�z���xĘxoxqDAbF�j��'P6_��l4k\�'Ա1��Ґ%&�I�Y:�� (,�'iICH�g�SPچ�!����q\S��Tw a\¢	���X�����*l��^��D}��n�_��d�ˈ���-��oo��9L���<5��]��:M���uS�| ķ��n������yO���x���P�s�:�H�INdJ��X�`�����֡qTat�q����o)]��C�� �!��Kͥ*U��Y�f�B��/˱�tm�����A�o:8�#n���%�n	�i|�� ,Z��p�׳����i��	�̬fp�i�o��`�>�:���w�K�wV
T@��[��=��9��L^T��I����O��d�S�a�[���xÁ9��'e��Zs�}GƑ��Q���~�<�ڙ�pB��C����Z�3G&�'�/ó�u)Y�A�7��}w���C:�,�A,}��i��ھ�l�%��b`*�Ȓ�c��'��J�?F E��r�H�eNz���ǥb�eO���m8�D��	�0\���?B�̈́��~w%�j��d���J�E�@���s��nΠ��!ua-�A��ں�#�~E�O/s��,��V��<>'5�<�rTar�x�)��b�6���^Y�_�L;��y�5�6�^%�E�"d�1�6
�b��9=�5���T�;Ȁ�F�-U��UJ�l�f��p����T�W� G�ֵ����%{�,t�w��������D�7���x`��tK����b��>o��]=y�$��_g�^_ډ
���o����j~�w�U3_D5xH���)o��P�#zP- ��u%2��ь\ ��
Yy�ȵF��U\��}�SV����k������ƌ�4��U���vN��2.��<���.��R�,�%����<�);i������3�R�b4��	��v[�3���ۿ�f.���]F�L��v�Oڰ�K=C�"�4:mQ�^-�Iy�JL�ey<b��D�b�g�Y;w��P.��6IޔBbh@��1�tij٘�,ĪC'�9�&�+�w���Yb�cG2���;h�+QM����a,�D�1-�~7^۟հ�M/9���)�^o\�O�<�r��]��$�Ptf]\�\E3+<�<J���t�~�6�)�Dxf̽�j��&|��qc���̊���1�$�3�u����x%O$�t���p��Q��T���l^-c��wC�6j@�F-��[tv�3-���~ZR>�z�RG��^�CS��
�6/�Z�^c;��^y'>/�Ն,��G�I������M�}Ia{���	�.�!�K�U���DX;|�cί��4�x�ǣ��:��9u%]�w]~�A��{J_v�t@���(36�TS�44Z�;=i�Tf4�A.xQInaS�B�ʌWJd<��.m֛lN���~|\�ʳ05���%t��V"�1&.�,ް���+aS��'1{���p��Y
�[Hud틲U�w��N!��th4�7p�(�YϠjE�8�����Q��Y��10�tOת��V�GA���chW�-=����Q�؛=8'�C�4�����������s��1��_�N��)��?䧼R�C �.A�3�Q�|역�c��@��	�Ơ��ۚК����E�<1�IA:PB,b�U 
�/$sh�Y�����^�v�m��r��eSؾ��5hq���Z���[����F��:ڇ�Ji
Y^piJ@n�j��3[2`��Z�}�X���v�@G��%��+:�)�:7�3�Q�v�t���pb<�(b-����k/�T��9I�P+�h�	��:(X�To	'dC�{�se)����IZ���6&�/+
M��ːc�~��p�ұd׳RYg�.��W��b��S�46<�/��m0���峇� �%�)�JH��G�fB	�+�W7m����nbM���1�{�(> �4,��$�Đ��M�tQ����pβ���Ҋd�#9�s�@4O	�#dqI�_p9)���.8n�`�B�6�ۗ9v8��ҡ�� �#*�YG���cR�vK>p���r󙉖�����,q5Q;�9;p,��X����Β�~`A'I�r�{�&��I��|����N������JM���ڦ���*Q���u�Z@��u��.tZ�������l��e\�ȴf��qS܊j��a���ف�,O^S%�^��4���jx�W�%��2�\��,���>Hq4rB�Η4�?�^C0�X�p<w�x�`21�v��]�ȆY�bH	%*b=��;I~���t �����P�/�Õ"��y�*D[�Ӡ~/��~�����
l3���h��IO]/XI�݁:�-|�����t�`c�ֹ��2�٭i�J�W�
d�W]��vT�����$��/�#�:�NP<{5wT�{���rz���Sjm�@�<a1ö�`�3���(��h~�����s��{�.E;y�m���d6�>\����v���M�4�R^ �GyH=P�)�4թZ�.�q�^jk���դJ
08-��l��=9���u���#+�N�Z��!l���:���T�y�ֱw�Im�5-4�1�t�Q����D��A[����������!�َ=[���/|�A:�S/9XT�� PJQǣ�B�遪�#�t�]�
"�Ă��[
����E�1
�zY�PDc6�\��8𝊀L��s��4޲����G��,a�{���oNJ���#��c�� ��R _-�.,�i
�����X��jH�m�����|��&C��� F�Kj��ɨ:lݑ���8l�2X��Z�mS�ݙG�R��ɬkʞ]�Ɠw3��b�i�ܖ�0
��	��y�9���HN��9	�`D���c� .�q,�͉�s���Nv�.�LR7��$5׍�Q#x���16���p��ը�1uS��R��/�?�VP�NBR|�R	��R��/������B��+��>0eo��S�ϸ��6�:�"��\V�����FL^K�
ZQ&� 7eS����Zk_��B#v{�۾��z��B�HLK|�}+ {[b�{K%��O�䖖w׳3�xٕ���(��baJ(����!�~��Z�WX��͂�� 'P�hG��Z�|A�S׍�P�4��q�,�tر���V�z�^�M��`��a�4e�����.hkA��X>+;/���jl"���g:H5qp��% �O�%�n����G�ro/����I`l�Rf�����Qi<9*EA)��)��1B*���Y�5�="�AZ� *Q �/?�7	`���LO���D�e�܆����,05C��m�IkIvm�cw��]u:>t0d#�w����@TC�uO����s��?�O?.H�Q�3����f��Ǣ�-	
mw��0Վ��!�RH�%�T��sJ�6v�0Z���c;���1X�V��i�q:~��ql��W��0���@�M��j�5�����.������"��wџ蒮�����1��e(�>��z�6���2�2��᝿��mwr�03�o)��R�_s�nф��wS��+�!�y��+fV^͔%Yp~�E����{�Ţ�"��4��_�Ԃ��_�,�y\J&�ݻЙr��e����褚"����j �fu$�ɋ�,��vK)�l��'x���dLnь��a�&�f�f�pB49&ؾF.N|�	}V��6z����dյyox�-p�8o��x[X�:���L��%�(�wi@��<m	��v,Bߟ����e֧��	�:A84�[x�|����A� ū� *�L����:��Â:��N@L��c��jp�����ŀ�|��ь�$�[�bgT�p������I�D��	�n�Ƹ��JT�Jy��a��z�m�:J;���Ҏ����!\��*��Rw��?p�#�]�q3�~���2��X��B�WTjTU�-i�'�gEC�D->���XK��=��HlԏM����S�.�]�/���(Z��V���U�$a5�I��ܾ��^\��4�/Z��?��	o�E�`eȖc���Wg߇����d��DhG��>{⢗�gs�.+mAo�q��oF�N��ysV��9�����2gݜ>��ɚq���p+�����x�}x��Q�wL�|$yx���I��R����@{|R���?�֩���8ReMo�(>���EK��[�s��y�:����'�5���.��P	UbT)'2.L���M/��o��>O"NPQ��iD*z\���Wc8Mf���JKw3o��򊙄�xB�r�����۔�/+Q�T�h�)y$a�>�Х+�?Z�c�I�:�h����Q!���֛>�L�1��pS�#����K1�����+ʕbF��tR���B[9͇�
VC�VI �yye"�5p��6R6����:��,�o�DI>�"�L��5a�'�ۈI; 7�b���_�a������IۑX�]+�"twزl�H���p|�h���T[ �,f}}�`�u�Dm\�J7-X�����p(�1[��҃h��3��o�f)�]f� %�3^r<���V�LB#��Y�ކp�Ə=W̤	�>��AT��]�-*��n���.��1��tҚ�<�WM/�z�*r�pfbIE�
*X�G�G��ϳ��I���|k��5n\��m&�T���(�xE(dyq
�s5ڭ����K��o0���݋c������4�F08��7R_��Z��S��xI!����g�ON@�Q;�ߔM���1A���]'�V� ���,w��R>� 7~�4=��cɊ��)��C�gY�ȸ�=zO~{\���+M&í���`���T�a43#� 5��M���;P>b"-���()M�>�� o��w�V��0��kG��kts��5�heS>������ �pB1n��!U��%t^�;�������)X"���y��������)��12~S��v�k�G"~3'���T����D0s����#��R��B�ҊP�	ӵ���r�v����!�Fp�o}j����5 $�AΚ��)�'jtUCG�4jR�1j��V,&_��i&����@����7����A���%)����`�;�n���2�t�,�%h!7��Z�ˇ=Bĥ���G�0���'`�������k_WƝ_����U'�vsr�8l�ٓ��ˮչV�/�� ��t�H?�FOߌ �P��M�5���k�)G�}�*�i{Q_;~/&������;�ܨ��5����H؅�d�';�i�	Ur���g,��e�,�:�{!��
@b|��|��5�PJ��.������_.�g�Dq��0�a�K�U�o�h���gQ�G�y�d�yOu�ն��d;��U^t��Jt�K�O�������ńe�r�u岹U ���З��-��72C\;hk�r�+��w�s��?��펽��x~]����l��0��X~��MN���,�bƑ�$]V/�~'���z�nX"��A�$@3d ���E�[%\wG�C$K�����s ä_]a2��j_�%���HÜH3��vI��4��UQi3+���&U���ൂ��UB~�=�S)(��ŷ�-K0gፒ�x�<��$=I	�Z,����l�;7��$����qճ[���~�U��p$��5W�R]����ܠ9�J���/�8���P���&�q^�;���t���ϥ�B�<�v�^\k��$�ft��r��l�MCz�E�w�ď��ᛋ����!�;�:�������,�N���Y^K�'��
-yM����j���"�@��G��0[X��^��&Ť6Z\v�% \c��lnt�a����KC�����$'�9���X��D3�t���|���w2�2���z�nc�$o�ۭ��=�,²Nן���?�)>�I���W����k�/tl&m����w��ZM�Aރ�bX�-��6�0+g�Q==�$f)�q ���	p�Q�e����do,�J�L���*Z��o(ޗif��LK���7NpZ���:뷼G�U�y%�zA�k��v������Fe��V�4�4(�Z��w�ZتT��ą��9�
˪����u�v���|RD:@��_Ar�����
���,���Ej֤g�x�$Pw�#����)�Y��h��͎R�,�ܯ{�3�)�O����E�y��R���gU%{����\�N\]��L�G3�_����"��9P���Ǭ����/n�B�[�a�	���R%&%g�o�{���3;��p����'�}ӳ�������(���|����c�
�@o��`�ŗa4u[���A����c��Q���V��@$MQ?SPH��'��}�>�]�����q�_f�HWG~�4�K��Bm�y�F�a0�j��Hr���C!��@(�T@�M�%K��EWm[�1!�&��/��7YT�_w�h��%��N�����i�I��$�$��bXjp�F�o������s}z3�?����`�oqW?�Ѳu�ɯ���|N�e���t{�,��n�	m�x�h�Ί���ز��}�~�q�� ]R��>p��:��hŖH�Ǯ*Y$���U٧L�[��G�j4)2�7V�"����.���:�@D�X,�h�k��_x}7������+s.���Դ*�����'�(v��� �t��.[DZ��$K���6
u��ۈK��/��K����[PC�p��l���a��Hu.��C͵:��##zZT,�L(�����,�d�-��%
�[�-
RN:����������-��qpɅl1��*��A�#�Թf��������,�I���&�+D�I����_@6��]h��8>�q&���B��r�ȏ�f��rm�a>�(�v�#��ը�U��C��$*D/��{�%z��Jpa2���ϩ2����-�������P%�0/���$B0�e�z��+�p�>��~>}���,�/r��s�����x=B�r�qj����U��C(�K�T����� UO����k�X���2����XWW5J��}͗d0�`�Ά��>R�`��Hj2IS�P�S]���$I���o�'�cB�>LW3�i�t`�f0��{���Er���C���lg�0��\0e�=�%u�.��硿�AH2�Ǚƿ��{[�,�Al���C[O��KL����dg��]���S:�����+�#_�/4�m�������U����i�vp�l���k��[*�����;�����#���k'�|�(u�1�5[�௴7��\�L�w0�Kx=��O0��$����`���kY�-�,���"Lq�2��C�\��:z-`��S�4[~$�g?b��J��q9J8/���d��6P`3��3�e�W�M��ՙ[�$���*`�W�7H	$��k����:'�2�Đ�P���c۳%v%lF�2�r�2���fyR���Z֓�)��˗-|�q�(
��̋L�8��̜�h?�Q�פ��<b����;����?ۋ�ǈ�j�aO�֨�н���~��o:�]�}O�e��Q��0�W�Cf��q{0�DQ��4��G(�nOĥ����������1��-E�������F���"d�n���/ ��r��82�}��#��� �9!M�N��Y9
Bb��������%��[<�*�C�3�<����ϣ�ET�57�OAz�I�W��5t�a���|���l���!�v�Q�OWK�.F��Z�z	8�<�� LY`$U�P>E^�kcS�D����2ɇfC��:��x,�t�*����I��M(]�a�/'mFk��7B������D�(*�U[�A-U��zھ8Լ���/�;.8U������L����(l����ؖi��J�y�:�����:߮S��B�QEd4�8�#��	Ʈ^�������b[�䲶<O;�Dj�k�	ɛ���ʏ��/�q�����M#�$
���H)|1��H>:Ww�ca�2�9�
b>f%�G���ֿ�D��d�}����(8�<�@NK����i���+DɄ	W�zǦ��c2�?����i�8���)���¸XK�ݑ-��ku��G ��&qBt`.Hy�]P^k�]�Fg�b�å��v4���3�Bu�wP��K�,.�义�rq��ˑ�W-Y�nG��t�$T���ն]gL��d���5{"bf}/����;�Nҵ�/���=����42�s,뗐�l*�cs�96��NU�i�~����F+6�l"����X���
V��/��4V�j�D3��j��.�Zf\h�d�v,��^�]��	�Κ�}L���q�V8��H���E��H��h??CGa�o�2YA�/[�4�_�"��i!�\=D��dt����`�g�������g!T��p=��.�N���Y�|��۳�C@2���>8�V�a*K�vo��$N��a�1��/��XIʧv�������u�6�	-8�`�5^�G�_��](^�����]���Z�h�_�����C^�LR����c��� C,*�2��p}�?�)�8�S�������������%�ĥ��K�e�`���+�x�v@ЫM��䡪�0~�:- 1j$=�����ي2�/̊�-�2bn�7%�5u��R�c�0��^rb����*|AoժV:�M���p���x��;��Mwf�Z�OR��;(!N1*m�.���Hww��+AXi�RY"b��Ts�L4�qμ���F�"�D*Ӎ�G�aU�)�7Пtv��c�M��7����9��9V��/����edn��`17R�^]%���פ2��a��o1���]oʧ��K��#.�f84ݯhV�B���%s3&s�wI�,󍃘����+C���ۈ$�z�z�7��o�A��bJ���6���k�߉pb?��Ѭ����+r�Յѳ'�h��בƊ�P�b�������S�@����Wu��rN$��W�M�7����1u-A��8-~L]��3[E��������+�n��6��&�O��X�A�^��S� �K #e,�{d�R)�A`w��3"w=wY�TK�ꢡ�vu�7�1�z�oiH&%V/�AŮ��-���JSP+p���硺2xCKC7�,��ό�S<E�b7/u/?����r�u��s��������.H��Q�g�ʪz�� �@ORT|"�;�؂�}f�!8%>r(��|�����|~?�H��Sr�[�c���_��	\�7~�T!0�w���K�V�zm�#J��.����P�J���B��?e��`6=��Rׄ�视_�i�+���9s ���-�%]�9�v�u����@~!7��+c\/bG�eb�����&�[α����\]���^���:�^ ��6�		D��\O�D��o���"b����N1<=7�����\֊��d�P�l9����ءD�u�a*X�U:��;$@�$�Πh��3��6,mK���7��9����N�N�x���yo��dL����(�����߈� �E��	� ���?�OV����A�?�]p+{,r����7����M���uwٸ��_��tF��6}�$�����ƓmJ�	��R���Ĺ���6V��F#�ن#�7/>�hp�
4ľ췌�%P�	c?Nn�Y��,�;�W���uP����d�~�0�PrH[{�����cG�<�NF
�;����U5�n�K�ى*��V�{��*jO�/j�j����C�:����l2�X�{�\h��;��3���
��Ų{Q�<g��Y�y7�TK��USs����4�|@b��Շa�>���,w���¿��_���A��h~��7�f��w�Ő�MV���S��t-�|��/'��L�5U0�O�ܐvo(�#�l����Ű��Hj���R�UwG(��=��CD��;�����5ތ���ӏ�V�0J6r��o��3��k�ڙ�2���v�	�i@9(�j� ���
�<c� �����*��N'7c<R�հ�+I��J����~v�����s���BlG�{b��2'(w���
P��t���c:b���B}�Y/�����'���~�B�K�;BCk�>>z���rjn�1S8v�ŭ�56�=2�:�mb"(���n�����%
����TfvXD�dZ:�><W� גϹh%�#��e�V*3��=����$�� 0��/r�^f#��)��[�`1�'P�%��m׶�PA�~�����p	����3:8Wb9��WԽ��|�
��-�q�2�Ժ�5W��]��;RLq����$���3uѷ2���j��#�-�W!)�p��2 R=�6��yo���I����X�Ko��H�(1MD�&�hj3�Z�h�'����a�$F���b�!osِ��GЅ�U��������U� ��C�k@����:��Iu\���:)Y��`�_7�;�3,,߲�����ыj**��"�"� �������<��G�äLaH9=o��v��{e�����Mׁ�,�-��wݷ��(����)*9mG�|���������#8�Y���EJm�m���� ��T��m�l�^��۰������q�}�Z�d d��(����Q����lyit�V"�Vpy��V�KpO�r$��tr�/��[��P�mI�yv��>���p��{���*P������5�gF"{���N|�e�tzP>ĥy�A����BQ�@����|V�����P�' 0�3���>
�f���UD�u���%��99��ᛷdׄ:F�Ҭ�����M�����N��|Õ/����̘�9��>�%d�,�]�!ה����kڌ�E������N9mK�~Ե��\G��;�f{H~#�'0�dU������T�GH%eD���B�J$�<������T��~l��W��/熳 1����k;Y,�
�j��.+�Y��7a-�D��6q�_����v�I �3z��>�)Y��+bDk��0�AE��ϋ@�10�S�</r�C�}�{%L�0��l/Ak%8h]�y����/|�t�6C�$��^�����2���)��=\��G�hFz�&�����Ȗ4`P&�D{
�p�����\{,���e���4{cC���������2�m������/�|�$!�i��+x����a����o��i�|��l����ꢶ��J�ƽ��?2�z��F�i.n_wS�-��.��])��=�[V�n�7q`��By���"o��R��n�pR���A宵#�	��~�]m봖�$��>�J*�����C��Ť���vIHPGg臲d�%�mBd����A%��:�q����]hU��~EKEF�&�j%���qyaF�`�{ˏSu
�/95�^�ј�V��m�=|SZ�aSf��=��w����R�� ��%��3���Z�j�&w�<�J�㗇��
vB����g�/|J" A2��h�.Lŝm�?������;��Q��v����%7&�
�l�����yA�>�XD7���(���
tY��'��©e�ˢ9�G�p#�o�f�'��y��{Au����p��\��(�&����O���)/�DK����3M��(2�@j���ݯw?�Ʋ\/�q��@�$ߋ ��w�rUm:�u�8����1\S7(�}-OGy-}L���&L�����P�L��M%�m{4u%����nö@��n|w��1��,'����r����Ge*���v�Gs����Bv�:�g�;C���2�>����%�-������]c�[xyi�^``Ȝ��]a��ZҐ��� �^�{���r7�+2�����aF^��z������f�c�B�̍(���{k���m;�َ$@D��9���:`aa�%z')�3^?��Q�fT�����a��e�T%v�ϿOL�Y�-$BE�ᠴ������)�H��n�
r���r��V�X�? F�E��ĝ���=�����WwLO�;���v����#�mճ�1{B28BK���Ơ�}od𱭾'��<x� �_��a�j�ɐ����D J�6������}������<��%�c5cXEq^I�}}�)�t�?CDߌ���.���l+b���R1���IK���е!/�S��hp����'=`f�@D�B�ν���Fb���=,u����M���;�Rh��+�v�H�>������ÐO������e����c舭c���å����d��y��J�*[��r���So:�l�a����m4�J,x,��-a�����"���7EEZ|��Az�UcE೗�u�+u%\W�o�<�G�XC����j�)Q���3S����-DQm�J1-���A�����% }���i_R߻Z��D'� �_
��'N� z�#�&��+L���ͭF�����)d��B��b	��2�}�'�[ɽ;���dl^��I x`qt8�wG���Sx��.w���q����	{R��CP�@-|&��K����Y� ӟ�����$'�3<��~��TZ����`@.�z���)��GbͲtĬ>�^4��jJBjduð�K�Y!�<&Š#0����%���}yA��Qd}�3�ܽ�`*�K��uj}z���t
����W���3c�̆���9ޮA�	ռ�xZ�����p^���yiL��Y��o�+M��\W~���"�iI��(�d��J@i�Rp΅��sS��	\�U����������I=��wD]"> �DZyxٴш��ȿ����B)֣?IZN�H�G{2
=����4�����>����"V!���:	W>̿�K���h�a_#�)�'�L���=���K Z5o#�W]vi�hY�]��}���Q��1�(��������,	�ﱺE¤�G�!BZcX����M��1q2�V�Rڂ�������Gob��o���X�	��%?�\�z�lhՓW�#���fq\m�h羧ԄC�2π]��f�G�?�G7��k���'!@��>���0��w�K���=�vo0��E�ؤ��s0��o�f<ԏ��bx������Yn� Ϙ'j��.���F�@�(�,�l���h��,a�М���ߵ����2�������)Tz�#z���"�����!�����%�Y>O�����Ư>dÙZ�u��ģ5�@��෹�e�@�B�Ru����o#E���D���K
�ڌu��S���
�������.	 pK^�k���p��t#����HhY��)��jf
��R�x�~�;R%:|�*���:i����w�L�nb��CK'�[�u�E�N=��*�-���T�#hEeb�.pz����T��a�(b����n�u���4G��E��S�H�G3u�,�"��
����E4���*c9�{<c葁�A˫�(�Kt[���|���lm�,���ݠ\�o~���)����A�atR?�1� k5i�OOl+�I�"�;f�=89[c��g|e�~��m������ӣ����m�� �U�CQ���d��!�;"�I� �V�H���~��}͈3�z�_�d��m2W,ɜ��;E�9ɮ�/������V��x4�e�����z4d�^Xh��/v���!��� L�s5<ΝҚ|%���R����#86(�.t�Q�g�791�*G�m��L��.F�Ry�y�B3<3��O���~�e.�j�3��e�	;�n;9ţs����0JÛA�1�yR��s PwbH���/)��VM
��Εrz��@�ʗ�(�q]yF���YjK�4Fg���'�>��Al�gfB;/�JM��Uwy���`�`�6�h�90�XPpؑ�ɋYM�R~�zGV��gn��=�� ����#,���~\?�P.�z���PCS��R*W�u��ʚ ��{�QjN(h�v/EGe��ߛ�k0VVY ��w4���˥�^_v�����GF�)4BCFƛL��uVcR����`���z�� \+g�� ��{d�cx<KB�u���5�[W�A՞;��C̀�/��d��\�/��Q�$5��.�o\%�k��QZ���@�ł\���Kj�q\��c��2�}MA�EY���Vu����q�ؒ��
�#+Z1�[&������4� a֌�;e�{]	l��:\���_4���ϩZ��l�����y�� �rҋ'Nh���S�B����QW��gʑ"GU={x��2�:௑<�x������$R��([�.�5Z���rd�t	1j�L���g@�j�c?��t�rϡ٤ �7	��'�.�萒�Pa$<�L�l5&,hā�C�l2M��zf� �,��a��6���]09�u���=g�I1?.�S��H�eO�5�H�l�	Y��׀Y��/	�s��xy88S��]�О�hI��1����'�$Aq���}e�����7�
��Ǉr��?1��N�s}X�8�Sq�ЁA��,�;zC��e2�#fI�zAf\�!�b�	�*p~�!�wE�����KD�V��mR��<(��-�t���(�"�S��L�?E'$y_4 �ؖ8��H����r��tKK{����cU�����?��ۛ���tg�{%z��;��?e[#�����\{���np�;���=*=)r䕊�'�۵XNT��L��w�t��:���y:���<�Cy;�)Eu��?g���4V6T�,�뛿0�����p�<�ě�i��g�AË%!���Ҵp��zKy*���Q c�c哰Ё%y���GӾGKc�y����9ߗ�'f6uu��� `�����Xg��4��^-�_h���=��Vy�&۩�:���n�7h�]�I�v\����+��r�cS퐽���?;Y����ʀW0���8_m%�v�ɤ���c�z��K٘WKI`n8	M)E�o��0/txHn����w2|���<l�?�Ǒ�S�{L*H��E�D,AJپ^�n�
zN����&;��o�rsзYӴK���x ��vӁ��K�룹6�T 5�\�i(qM���s8=Y�e�+�א7�����C5%����j�!����?F�G�s�}�j!�fĸq���W��S���-�*=5����Q��_�r��~�io�LV����I�8�����z�1W���T$FQ�c�3
���̄�{��(��	!?�������X�D#���p�!����'�����9���Q Y\Y�:��_�o�m������	��)Yy�'��1��V�]~w=��1
9L�z���i>��@ �k`1b��6�2_���^��.UP)Z��OH���:.%��UJ2klⶸ��q��$ĕl���dh���X}&0]����ȁfq�2��(x	Wr1t
��5���U�ˉ�D|'$�L��҅陵!�O�;X����n����5Z���x��z�J�}r�����tM6g����|!�[�"Đ%!�Q�k���A�L��/�h��1���F]���I�cs�
�P�)�=l@�X*�����	���;ԍ#�Fu;Gx�;�ij�w��Rs�&�c&�)V���aս�� �屑��<{ ����i��S��R*�F�`~_���l���2m �x$k�9d��mW[ʀ�G��c�����O�`�,���;8բl.;��]�V+��z̋�_�cW�����{U�-E���o�#osx���cWD��[92d���{�m�MT���l�Q��w2���$���-�����g���{�Tx���R3?א��/,��Kk���;��
"�����X���Nd�j�.�-<�{�x��.}S?Y�����ި���^<dx�f�l�=��$*��C��I���(���&5��_�=�W�L�V�pؤh��:ts7�U�7�-�?�����V�z?�n��v7�����(ܜ�����"�
��,9~g�[T�9 x]�Cw+�ݺ���E`w&
<�-�M��P5C��R� h�\P��Tq��ҁ�_ �J��:w�l�=d�O��,�K���Д^��HrR�����>��lƄ��U�Lf�P���5̯JB7L��#+|Ӯ�ч2�HȄ�/K_:+n$�ȭV�F+^~E� �U�t�@�U����n�"���#�e���]*#փRBU����5�*������c�wZ�sx'�e�
M��.������K�T/v�K�&��~l0j!���(Z/E	GK�B{6*���0k7D�9%�T��,m�`��S,��=�S�e�|k��rd�Cfso������7X�~r]X��{�I�'0�nm��ˣGDȁ�q�t�{���Z��$�����vF�� � :	��I�2��06XN��!�7��M�sd aN@�����e�Wb��5������`!7�]��N�?�$L�j�B����!�Xؐ7Q�X��k)�d=�����@̜���W�qLވ���X"�q��g��փ�$��I8�C?$0��L����M�ɑbƵׅ��2�:�s����X%/�|i��J�'�����F���`�,��u�M�1\ �K��	|��&����庝����Ans��X�%��	�5�1�ގ��_8�u�'�7�t�<cv�=gƯ���mVior�6�O�I&G��0i��
$`�e1�`�f��79��".KN�PM�G1�M�k���oq�FX������%M��p�[��x�o���_�8���F���������.ų9xO����MN��_�՜�Q��\o��Gxu��g9��[��c%��J��q���!֚[��N��{D��O<BjѨ�0���3}L�jX9�G{M��H��}��T?�4:z�,?�}�:]�'ԡ̅�%�GS�6� ذ�d�:�n"1~��I5�V�u��G�y_�J�r&�#���pf���y���X���+i��7�J^@q˚�������U���
ZR'����6V����W���|�ӱ-+�
LeYY�t|���D�Tj������*V�R�I]T�6���������P^BZ�x8�w��ѡ�a~�U�͑��k��T]'Oj@er=�20Z����Ƿ���P��Xq?a��PĠ�I�����!��%؇�������'���k�b��EҴ{'?茐��;���Lp2���B�+%�Ӱ�M��1�G��xK�!Ρ8Q6��LVF�<����1��r:�rj�9[Q�A'����TS��/U����W`��G~��|�0h	�c.)���#
4`E�b�s����Խl����L^��5A�ʀ坙Mm�__��G
X��]sWmKB��kp�Es�+=U���G�[�;��S�%ø\l�3����*ab������zn�W�u.~�Z����:B��Q�#n�P��c+�M��֗G�ָZsE�`�QX�fK�s_V��%L�༤I� '�ԁU�B�B6�� �i����n�	�Tb
�Σ�dF�F(��` ��F��A%�𵬶^��AӔT'Ί�L�I�镉��C�bs��@��(R���CD�R� �7$j9iO��:����EzyG���5��L�!e-ǟ�{_�� N?N#��H�	G���bq3�WnX�x�q9:~;w��
�V���J	�3�ЈEd�\���j.����	�}?]�y��A�j
d+����i^A<ϫX�,�=r��:�4����l��~i���H�8j�=�VM/6p`��X���Z��eS� }���O�X*}��+���+n�|����K�:�@�����b��|�Ht;Xo��ezh��=�-�D�g7��uz��A2{�V�l�+_QɆ@�Fa_�(�_���I����Ũ��P��1v#Uz��w(|�8�{��0#�D��Nu��.��rzT������ pF3�\$�	|����F�6� 5"^v֛m[{A/������޾�C�����Ho�u<;��y��h(}�C���M��d�Y���:�^�gX�2�v�4�����h=�;��	/���2�5Ĩ@eXI�Z1��z՜�7�Lo�� �!�K�t��oh�{��O��M���`J��:�!�_u�{��}�g]{u=t��+�ɩ�T;�x�VX�O����τN�t]��~�}�Ǉ�ڞɺ�r4ٳ�\ÜH߯P����E���4?8�<��uYa%{��+U3��@>�ٕ�#2����2��OA�w�~��3��g�?{c��c`���V��f<Tb]�6�$�Zll������2��ْM��k�Q�y�}���R����`�.%�;7��WFcd���*�j�:>��-R}q����ml+��Ӕ1Q����q��Q�V �S�%
�[��q��Ҝ�n��➚���SZ���5�<�����q�����?�SaA�Di_AhU�����}I�_P,�9>6��kʵ-��|wf��rؿ�&�n�(i�	���~G��q���3�%&��%i]N������ ��l"��#���6��󄾳�^�^�M�'"^�Nl���a����@�g����*����/��1m����|h�o��}E�����0��}-k�d�|��٠��M1�����h����,u~1���r̽#u7J�SQ���aH��|�T�85�� 7R{m��c�X1&LG�:�[X�7i'�^/�������W��⳩!q}����c�8����[�[�W� 9��	��gj�"���))�]��4{f��/�G�\���󗥢uV�X��ƹ����>�^h �zb���?|90���/f��"�y]`�4pe��<m)wF��p�X�*i��ۙ|EIo����������H�܇髅B}s7�F�
L]Wz� M���L��ݾ��[�h���K)�[G۾Ϗ�3^�����9?X)D
�K�G������RC���G/��Y�eX��s��(�������~��'���R6LC�wϪ�_��o*���KN|'�8�L�(6WeKhm�[�]������= 3y����v��m
F�<�Hu�.��<`'�/�
��{#1\�0��R�����iqi�P�F���y�X �_����o8y��]�A����~' ��u�����۬!�u�k�%���{y�<�ಷ�����.= ����mݲP��K�|��'^#exA���	��4�bW�Du��K=0 ���)X��i�~tf		��_R`�(/Hg��5�[[:�5��x�_�)�jƔ�����5�k4��OR�MJySz�E�=�l�?��ힻ�7���ǡ�=�։]p( K� 5�K�H��n�2�R�UAur
O���	t�O�-?��3;|\�#k��w/S��p�pb)Pn3(��k�P�1K%4Ld���,E��<lv�u����8E�! �2��)ߊXd�o�:�1	qM��S�Cӛ�D���]�"6�t��#�x1��=���hMb�?�̝�c���AŔsI�`����x����ݍ�X�,چ��	�\T+�1��gly+8��|v9{5
Yq D3���U���"A�Ion>�S���¹^�tT���ى��C�g#��uB+{�K�=�if��)��)XtVtD߫��/�S�tY	X¯;i({�5H@N5љӿ$)\ ��JJH��x�+��;�Q�)�΃*n�aK�	��p��+۬εX7_�w��E�T]���o���5��X5��^��xH8�%~��WP8Oj�5R��3���^��ޭΘ�>�U�q6��ܘ���������F��x%$���l�AP�f��#+<�#W��+�
Kq���AS��ր������DR9xe��/�%��g��m2�>i\���s��ܢ�_�^��ơ,���;؛�/�1n�f< �<�Tq4S��t���v�R�����&���.����~��yM3F<obUC�2(B\���÷�ҌA�9&�;k 3
+h�&���ܸ���Xc�JC2�$K6�
��^E-�	�pyMIj�nG�Q�e��`2�)�����(_���ʕ~K'^ +�'��
��X�A��vS��"s0¬�i��Q,@�Rӿ���I Dŋ%0�x��̽������6��m��v��}ت��k*8�t����J���0� I��<�L��[�gm��NF�\G�Z�"��H��//2��VNf���f�� >���O���O�#��)� U�����yN�fw��Y�+Xf�1X4�gJ51�S��~P�~�O��m�FX�´�o<�'#�����?(<��rݳ��2ҧ*.����׸X������g��HcO2)�@	Pop�ޒϙ��&�*�����R)�;�Ξ2�U�� 3���Wi���%�o����)'rt���9�wx����)�a[E��P�Ah���p�-�[/�N;�G�F������+��jv�fF�%�	���t䘓����I���"a�Stt�1	/�I�?Z.�*��v껞�hvĦ1/���]?��ܬ6ReT�(bA�K�Y�����`��z� �3~��W��;]�3�쓮5*��8��������\\*�rE·vk�ɃW�L��������\G�oX�rd�-�fL��xc ���Ԙ\!�RRe����a��'��bG��f","���<���QIS��ȏ�u���ʬ^�!��H����ݥ�/��1��G��nT��/��Et�$P=��{CDؾE�{�����#�*I3��r�ïm2���N�?FRBHN�V#�A��	��q����2A����?6ᡙ�O���!P)Y�y-%��������Ay
1l�!r����H���H�v�IG���=����:��it���.�ܬl���ӊ���c�1R.�f��՝�=@�ӡm������f��O�B��e��!g�k�k�|y��Y�	�DG�m7�>]@r>M��"NC���u����8!�o�nV;� Y���D$��b�r�Os��: {a��NK��q���f0��/s���ͣn>\���^PVq!���u=�k{�&�C�x���E�����4�Ic"-��L�`��/���������n�#�}��j��+{����nL�4U���v�H ��	�$����:|�T�w�A���-��K[d��B�ʭ&�ˇ�O���R+�S�r�����Ѳ��V���}�I�R1��m�` ��L����:���aĩ�y��D�_���Q��[��}�m0�S�r:�Ki�����Zz��>l��v�κ[S᳅�/�8B���J��l��(�b�қ�� ��v5���R h]ܝ9����M"+���1�b�A$6g���`��Fz�������Z���.b��$�b���Fe���Ш�Y%_�Tb�:��w!h>JO'wg��?�{�n������H����ĔEɟ1��Ǌ�;mb��z=�������8�D�����D:��#Rv'���m�V�Tr)�NxKl�\GY9>4�nKB�Ƞ��x/	�߲���Q�C�2�c%�i0�7�Z#� �ѿwQ��&7|��u�y����Asû%�х�E2�*
[x��C��$kC�d����?��d�!�� �:�4%���R��s�`bj�V+[*�f�y��]�}7y�ټ�g�EZA��c+���I�~e
�����"f�o�Od�j�𳿹n��n�|
�#�
i��
v���f�_K?Ȁ���H߭�=A�zx+}·j�l��!2�p �WO�Gr��J��^��;)x$Kܛ���1�Yy�g��C�������H�ZAeO��0
��xa p`�L�ѭWv�mH��$ً)-� b�o9g��Ag������N�"�M�(=O� cq�5*�~.3��_����9�jܖT��d����+p�j��&��L�еQ(c+j�-���l�M9��F	���=X�i�'!��4d��6��U���"���5C�0��\x��)�x�dN#����Ο�h�T`2�ʣ�g9��^�ٰ1�G��C�j�iyڴʪq�Ppy�v��]4��[�h2���ǳ�w����b]tEV���/���C���[gu���nzX�?�PU��l.��S�j2��vd�f��'�P�� a i������WO4�u��ٰ�z7cݳM�8۔9�����b�����3r�I�/�C�����G�9v���äj�w{����臂�Lݵ#�:<jl)�EDӾ0KU	'��ok�w�H'�vN2�����IxZ�X#{�gyiu�{H[	�æ0�V�0��@��d��83(kys��_N<�/�͇ڭ����	oq�E0�1	�`6����t;����7̀
�)�p��,��u�Fe��� �f��N��[���9��泶G�95�ɡs�KG\Bf��YN����2r(/R r��GL�ƴ\�#�m��k��k�NY�֫X�s�3���:=u<���� b��8gj�#S�jZe�*I��Eh_T����	[� ̒������r�v:D�:i
�;�U��S�k�����gY�2O��b&�0�z�'p��@|�o o�����죄��t�<	�|b�e�>Z�I�f㑀�g
�m�虒I���s�*
��U�X��X�L�h�Ҙ3��\�'�(~��Mk�c�����Ga���@�(L�N��L�����HzFHh��`�1�5b�X�܋9�ee����0H#^զ3'�	񯯪*�>���9��5��?� �v�Ek7o��P@<�7�"tx«V��X(D�G���6�m�,ԕ<�����B���u�4���D�
���-h�Eڍ��$��Yȑz)w����eg���!9�?6��>�[T�T�����6 ���b*��o$�KB9�{��6������Z��ⷐ�}�sO��pl<���^���B�~TO{E1�H˔�ͺ�c��M�������H����O"m��y����S�7a��6�\O�c���&B��c�R��gտ�X�Uۺ6"[��A�Q�N��SSu�$�P��'�,�����ʣC%�-s΀�5"�ե&��f��}��߉|�����V-���\l
�B ��0��>�ц��"�R|�
�uj��8�Sp��:�.��:�q�Ace���}���s���ejq��<<:rEŁ�>��H��X��4�����
����c�`)�V�������v3��kM?>Z��[v�e V_ڂໄF=�26e
>(�$�N��WCP*�w���C���s򠷹$�1M��{��˂�ݼ4���T��W����F����佒u�Cà|��m��ըbGۗ���� !6KS=k��-)����g��a�~����t/���+ۅ=A�s���"���j`.�<�Ac0�,^B���녓�t��6���w�{�����[@/fFƫ"���[b"\iT�n�V1�R��0j�oq!��;��D�Uh�$T��d���'Os������%M}$
�)���|�c�m�����=�����n�pKPN�p7N��N���Z�D���)S`8��tO&N��"q����wu�0Q_,xl�'��`[� @��T�l ܽ�Q�E~�@�CP�吏�AX��e0���Z�qs�f�5<
�����U���5��y-¿����#�ϰ�����h�H�8ieG�|�9�c�����?�e ��wfM�Xoh�d���kejwJO�O�FZɲ?�9��
0(��z��@���.�E����E���L&a^�D�GNE�,{��]�Q$��o�r�ۻ�%6'�87��`��h9���AѠ��O�U��hY�m5�����=V(Ri9�߷E���`l�����!T-���j
�۟��} >���}��bd��4��j<����ᜦ�	�3K�%JTy&�a�>Wz�!��M���=�^�ʫs(�����M+|��Q$o��++��ԍ��W�����U�Cn^�y�}P�?T�|Q�,
Ǖ]��l�=�~u�[�!���4��g��Å�'�3g�'����a��a�l�̠鋀�}y`h��-a�O�^��#�S��d\'[��5�1Q��>���/�D~T0�R�}SҦ�R����z>��am�2t�{�7�aX������t�V����a h^`Y�˓1��RFYU*��2[�+�����'����u {N冃A��u�*(�3�wo,��)8w�`�B��p(��X��A!���q�'�ʅ���	������U�t�E�(l��x9}[y���!�=O�qG}o5@x*�8Ñ�h��F�Ê&+���2_!T�����Y�q��&��n3�6Y.�� �{�Ʀc:M�Wml�a�� ��;H*3�8��T/`��G�Ƅ	�[֯���8���h�j���_w*�i[���YB�r(�<��#��/%��ȓ�KzGo�Ki��W��V�����2�x�%y�|K#�W��{�?/��u�dJ�9�\Op�;lVໃ�y��,-Q/�d�r8N��_��6!
g���'Q�"��Nw���zcjCS��T��aTT�	�3��O�_#����#�z]`��R����$�u������C�]��+z���'�Qբ�,u�H�dzL%��9=�_��>��Ŗh5����6�6�}>��$�Tψ�VI��f�Ʉ�d��%��I�!�ڟkJ�91;x�{a����1���rl�C?�-?�z�-7��S�T��G6"s 
� V��|
j�+hʅ��8���a6/0R�:	˴�*Ψ��xq��fI�#�|� ���A�4�os��_�3g3�_�8��B&C!Z592G7�L�ڝ�?��r�q��ߒ�-cӓ�OYu��R��i@��?�]�h<|p�P'�*��:K�Ƴ��aQ�u�4 ��=kC�����`�I�qO��4�/��ϳc��$:I��y��"���(G������ݏ��+��E<s}>�9,K0���r��Q�LZN�	���夊o\��_�n��c�� �8�ܷ|�R�^�̭B.<�'%5���Y]z���{X�?plG?�1���*�A��/��d�,����C,Z2n��X7#^��k�W�05i�A=gs��\��
�T���0��f��bTnz�d�tP_d��h�߹�)%��SW�tt�,�"e�6�M��Յ���ڒe̵�`�%q�ڍp���Aop� &��Ԟ/wQQ�q��P%p���s���RC�n��(�1�ηZ�"�OG�.뾠����4��B =�gV�]i�t���P��Ǡ[�9���,X��)M,�Z�� /�؇b�1���\}Fq��w�̱>�cu�l!���xV2�T��&r���VL�=��HeW�)?�����"�|ޤ��oT=��(Kǹ� 6���1z���2�߲���w��a���"����<�h�Z�#�&g�m�< �}CJ���1s���^97�o�fzH�-r*H�G�M�W� �]����b>�Rڥ���X	�XJ����L8�)f��㛲P�p���Ә�i�]��Wn�����:�{��h�h)��ב|9ڸ�L��O�c`�-�h�u��3>��Mv�S� j�Qp��!���[<�p�kݿ��%��[���(_&����
�C�c�	�}<n�ـp*�v��������N��U��)���?0�>t��M$��HD�c|��(+e4������DV���L�]|��ۖ��OK��D�pDN�f��T����p�B���	5f��:HL��O�q��	mHsuE�\Ix��I�>AA��7Y��xx·��g�X�Gc��LK���m������V7x����$ង�Ïj�#����W�U'��r�T��_�K���'Q�6��=+�U�:�2�?�m��<6xB�3آ���CՁ=\�>�����zЧ��EuY�bQsQ��C̑�vUNx匹eDt�T�F`��Z �p_� J�'*��� %���F���5��s��C�����ߤ��=�Z�y���.��=*��(Y\�(��(o�0�3C��(z�zBYduV2��G��l��k����|*�f�S�"O��|=T�F�{���f�� 2�L�F���8��
�.��f<�<T0{��WD�1R���7À���#})>�!�y��u���
r���ƨvK�#�*�p����m�GD�bB�d�5!��RT��������/��أf4�tr>���>0��t�.��jP�L��^U��%&�z[�MY�^2(�L	7�)G �tџ�e�S�ڏ������#��B�V0a01{�J)�s�[F�Tb��Z���)����S��6Hr�[���,�-u�N+��f#8��8���*dSh/ٍ�]^�� ����B���[V�	z����)�0
��Zt����n9�ᆨ� �?���3V,��a������9�c.V�9����s�����b��]�I?��p����Ӂ�<����L����?��s N3C�^P�6�[h	�ܪ �˝@j��}�D�NR*n�}�73�Vau�
V�g�ۆ?d��V�L���O�8��^4��ͱ� �x"�]�Y�d��}����Ќ�@��O7b���"Q1��80n�`b�)d�Zuf�-ț[�h����;�;��Ç��y��9<�DH�N�˔,ab���'����郥�]�9
BD�H\�h�~�?"�`�h�*�n֊?Q��p3���J�Gi]� B��Q��s���f�m!X�Ԑ�����\��0ިw�ύ���TD�ijZa���0�Z!�O�f�^k�@��K�҂H�A�G5rE9OI�B�?M��M���8N�s�ҷ��v��ņ�-	I������J��F�R���T�߾�_L"a(a��1�+S<�ΡP�7"�;�J�;�#�Tc��Ư�G9���b�Wk�u3(�ѹoŭ��QY�<��!�_�&k��e8z12���ۥREYG�d�`Yr�K'o0���'�3��yx���<F��+;����D�t���&	A�9L���B�J�@�I#�>��LL�L�_kut�� Tԟ!^k�Z�`?3�tD>�O+��8M�^��Cwy�����A���lgx��ɶZ����������������^����dо�!�
��qÙ۠s�-�P��H
VCҵQze����x�U��S���Py�h+��D�!:J�7<�
á/����Jx2׮�ylP�QR� �@�R����if��'�a�*M�/��
�È�~t�1��H�:�#5b�+P��q�=%T�y�~K����>�7��m���R�qm
�����}�q��ҧ��(�m���/�̃J��O�.�d�'�ѧ8j��\� 1z.�}�q��6�|��o��P{3X0�[ЖωQ0����Y�`�3���ҝ���d�L9�����슊~�����F�f�3U+�D�2�5ʽtj�s.�>�i��hs���}R����yzLh��Wj�w�u�Y 'h�e̵A�gݡ`Vl#�L\SY���9!h�7�@f�vZ���E�r�0�����&�p,�T�A�~M���"H�����;�<�ܨMG���B�+��2U!�ҟ@���m� w��`t逐<��	F~�^�����l���u�&;��q��a(��Fϵ�*�#�&��c��]m[)��z3�x_i����-���@��j!�����;�y�TJ�g�[�c�`p��͢�C�-EE�aл�)�+vn��'��$�l�)6%Nh��W�fڐk�5ƫ��5\ô��7�g����%���1�d�χF�p�Q{�je~�ƨY�?��7�:��]��%�|LN.!�V]�IO3�sC��)��x_ Rް�N�"^!q_Wrb4s��5�}=�s#S�K���'�{u�[�v56חdV�jɗN�@�ч<�� �n+�čb����1������ݡ3\���a3�X��,�BY��'\��/T������LRo�ʹP���-��m�������Y��'�W�;N�W1��GH	��bs���S���\x�s4�1�����t�[���[�NV��i��Ƌ�Ϩ���dw�j!�P��m�v�9�
����t�2q-D��T��H�xy��q��=���~{	�,o��g⇞�"L�rg��vE�T~$^���6�xb�..�]�<,��S<�����6�{*����|<�Y� Y���c���'�Xht��K��bE��sX]�_;F��تl�x��}�d����7�w0��Rp���D��o&�~�ۑڿ�Hud��4�B1�$9�U����mh��$�J_G5(e#��fz(�"*B3�v@��uw�S
�ƴ�A��I� ���=��7���|��nB�t���z�d��6he���@t��3Q�;��6��2��� ��*SF�蓛��r ��I���:	L���6��&t���-s��aſ�>�sr^G�w�c�>N�<qP� zg���}m��5k�r��˟7�3�k�Z�?�<�H�B0Ĩ�M��!�3�4Q�Ms!a�eS�_L�����(��Y�?�����얶W'�S��8{��0ۜ�e��{z��ED���ЍÖ�5���/�u�� Ee䁥��a_���g�ݲ�����ٸ�!�,�`��X2:�'ll�at@�M�>�4��k��) !F�����~h4,��LNzn��v�x��<�V�4f%�f+[;�Y��n��!�57l6�v[}\�`7��w��������ݧv�s=�JU\��qd����A�IGd�����vk�(>�� A!�W�g���� վ�Gn��h}�Nە��ީ����DpN`���2����M݄s4��y!8�=Rv^t��H�a/�4�w G	R�e]z���j�����ӿ�e�r�8��C���Ӣ'u�x�&??�f�,��^��2(Ǔ5K�)��}��a+����	(8�w�ڝ5��v��ӯ����r�n���5���C�<�Y��}�S�kU���Y���PgƳ \]A
���݈����J�S�:�E�T�?1�V�,�oP?��۪�<��;�W,�;�WǑ�Hj�G왩W��o�����K�oI�p (�dʠeC���.�~}6���b�}V,��M�ʸ���hX��{S(�m���^T7}���e�̲�t��&�ݓl�# 2��
|��
�n&�j?k9����l�k@��-��OZ�wk�s�%�Uڙ> H�+��3U2z��C��g��+�'��LF��ٿwW�ͮ�G�9]/�"ُ��d�r�G|&�|�t�G�G������Pbp2�"o�9\�B��a�/#S] !���F��̋��L���a �,"�cfXH_3���p��T�/��(���.&�j���ё�oTn�ji��#4� 2n�X��(ܱyYu��N�%qZ��W�Ի,x^R}��w�`?o��*��/�
c�W�Ruc�?�����ةcK~H2����벯�ڿ�uZ\<��E����#\��c�-]�<5�8w��E/$�șӸ��l�c3r�I�D�B$�*�}*�L����a���I������慮�&�qZ��1�C����Lf��d��r��^�5�r�[�~���W���vB֐�[~�`���6��F��a�bqX�*%�k�؋|�V�k��>3`�]oR��PO�ЈS(�u~p�������&�����f=$VE��(U+n�h��u�6<Z���6�/���	�3��6DX�.lۀ�b��mP�I�	���n�[�v3���#^\��^=�����Q������*�C��c}twv0|�3�>���mU�/F"wJ��SK��u��❦������	-p�T3��e�c�!�a.����i���$0�Y�+�=c|/ʠ�cv�|���E��y��Ԣ�F ����ݦ}�X���ԧ呶���(�7M�@alk�S�?���5;�[d��E� 'p��ar-{\� a v�1����}�i�(I�l�J��.�� j��F���n��?�B4�r09.��+վW,�W ct�[HX�͎�N�ˉ�j� �Ä�V�oL�֟�ra��z+k�q+�R���,�I��6�A��7	�k�����mwl����Y�%p��3�q�c2�ܙI�/i��Ե}Ө� ����� \t������^�d����y�0���kZ^^�@=�xd�>�i�+Y�z�w�]mˠZѺ�4�J���2R�u����pI��{A�eG/��P�D�Y~wI2�����J���%�&?������u��9��D�{�����JT���Ϊ`V��i����i�4u^XJ��VT^Ml���ݾ&�2�j���'w���CN���2&�Ѻ� O��ecNIF��B�-I�\-����Y�ZaQ10�?���t�*$���r�����A�@1һH�٬x����=?��#�a<\05�^��@AH��P~K����7��ELk�7b�os�9�h�G�����V��[�G�|�]�4�����$X`<�̴�q]ڏH�+wc8����}�6���Ov�t�L��WW��5W���
ǋ����6c
c�����~�ۓb#��
�?a��ϣ�z"Tf��-gƒg\D�C�e(��ҕ+��R�X�O��y:�%-�4.{�l:D��r�_8�hy�����>���.��A���P$�7{���44@��ǿX4�
���uo}���@�̟����E����N3zh(ذh16���I��5¸��R~pv(<{[|S8Ttw��F)u�b,Rˏ_�?ɯ
t/韰��~.�(��k&�Q@�.�y�IҔ����|��I�~��U���	Pk' �G�c`a����N3n5�0�$��������Y+��k=�C�������;v� %A��s��~//�qgnk�wr�f|Rldw�ѻwܺS�9'���E{k�,��x��Z�������=���6N��8Om�����$��@��R�g٩��O��� �	̈��o��c����#�B�5��L<��5�`��o��Q�N��T��u�X�*���[�ڦp�f�8�"	�:K��9a[���-Yrw@�6ƈ"�^� ��4�0L7�d�m�.���̲��e�~���@�m�Gۗ�Ѯ�5c�C)=H����9��T��d"��=���H��En�q��K�Y�3/��d��KT�m�4�ˊ���� ���� jrC�^�2K��(��-�cc����#)h�=x�4\Z�p�(p�yR�X��6S�|�*4j!]��RA���W��p�#���Pj���VB�"T��ǥK�(��~�P\����s]�����I	���ʠ��A�x����~)~���	x�����f*��S���O�w(+/.e59KS�|�����;�IF�o/,m߾�i� �=\��i��J2�%m��ٞ�8�_7Q���&�'���U���b�ڪ�����!���ܵ��$�T�[?��h���FQ�@��G3Ѷ75 a����.��2<�>*�[c���F�.��
>-h>���ύj�GO�e?�f:�`��J�$��_�=�!�N~��L�����A)�6��ј~��B�@��O�A�ְ6�Wߖ�{S��k�⛸���OV���RG�aUn)��=N`��4�ê5(sWp�W�9����L�v)����K���j�\'��&�:܃C�Y�[��������~" L�����f��#�G+���]�]���i�p�(���\�/z+��J�J���`�ET]�y��mݮ�A�l!:�(V�&T����s	3u�֪�5[�~b͎6
��&�� ��ޡ��6����f��� T��R!��ee�JI֝�e��\�%�~��'j�}DAir�50���j#�Ny3���c�qn/rB/96,E�:H`�6w�"r���֋���kv��i� �VCI#o���r�)��%�99x-��:d¸JҢzq�ɻ�3M����`P�̖H�x*���7g���<�@�r����8k����"�c�'H��Ɗ=}�1���d�k[⏈1i�&��~� �we}.���r�Z4��5�O�#�8����ƑAz+j�D�w����%��6ԕv�sn�B~Eù�B'!??��*G��>3�.��}��a�Y�v�򾿀��K�� �m�mT�����|�~B���g�� m�2ͧ�O�<��2�GM39H�����Ebr�s�D��NX_��6�m�f�<�rъ�d]h�c��đ�!""er��}F5�ģ�h(�h��%�躭�JR>;Pty�ת���'����w�M ���D�x렼�j�n������Ii����Iz���rd��b�]�Q4���x�ggd�����5M'�E�ʭN����*=�z��W��5Qk��2Լ�1ǘS'Q��|��剙g~��c����Q��#8�W�^���Btq�p:O�k=�w!F��0��r]�A�|f��ʨ�������܎ȿ�p'Ǫ69ֺ6��h�(��ݕ��e�w��Q f���\�:�4N�-�`Ӆ�˟m�+��d����D�7(L{�����?B���.~$�]���ē�~���<�ΰg�hDd]Q�BXd��v{���KR2h�w5Z��ӣ����Y� 6&"P�W\�����~��mD:���[���C]��T.�ǋ2*-�pd�n)��_�J��&�Etׂ!УR{~��B�KW*Ӝ$�7��`9���y����J|�6���_��Y"�g�BF�&bꠈ$��F��LxAM��
�)M�k\®��ĕ]j�2��Rp
���̿B�M{F])�N�J�	��}���˝|�t��+@��͂��վ�a�H>D7�S�a�xE�5'6�po�8Ne��J��_�7��tR���(Sy��rD�h-�\��w�ݞJ罏���p �{�_w�@�!�>e�l�hX-��,M�[\X�_4VA͆,y�K�ܽڂ8E�Fճ�E�S.)�ѥ+뱰�������7V)&D����jVV_	�i>5fm	1O�c������0�w��!c��υ��w�^��Tem{0g����&�,���ǵ��uhK{'ǅ+Ań�ΤhB�a��������54\��[���v�̞0�[@������53݅F�y�J�MM����K�����o�������D����t8����+���~�~����yI����7G��l�)a�?��9��U��e��c$I6��� q�r��$���m�5r@#��|����R��.�$�i��Vƙx��N q�4��6�o�čj�,����<[N�4��XgL����߽�b�)X���2� �\�T�W[>���69��4���$�(ӻ�l�gzcF�J�Zt��6�]���*�6�б�ǋ�v���w���^��; ���Q?��9lϫ�!R��' �lC���H�0V�ɟk���Y
x=��AɎ%D�,����Z�پ4���n��|�w�Մѵ5��b?���r�R��s˲�M�I*�Y[�f�흿�����
���a�� ������tm|F|JH;3��1���an3Fl]�&/ܣu~R��t��N|O}i��w48���{�^%��aZ��(y�aqT�^bg+�<{V�o�\�� ���p��V�x���8�ԆZȖ�e=���uUf>U�G�D��7U:�$�Po�I\����z�J�.���0̘Q�G{��b*���� �)�8�6N��׭3G�.���3Z�n�	��'!丳�k�f���#,M���/�y��嬕�{S7|�j~��m�Ϸ��k�{�D�EdX�=cj�S����2�őY�n|�M�\��D���e�r���fn��8/��[��\&��r�7�e���ם����J
h���(X�0P!�)n��	��#��0��&��fp��+p.��փ�����B��[�-�j�
��Ж2a���$����ˡ���Uze E�.�#�k��2x�μg���{w#~mq+S*B��e�[V��9�w�s�����qM���ܬԎ��]M�S�'4�)�J?���$"�����X��yeb���;��u���q��3sk�<dK�lmb/	��gY)ᄫw�A��{�=6��E{��2���3-c�O���~<%T�~X2��mn�r*˜%�d�������Zv�k��� b���<�#��!�CoC2���v���E�d�ٌ��R4y�K���4��]-�e��H��	[j^8���a�N�XqT=r
����~�1��<8"z��wU�5.�]n\t���Cય�!ʥ1�����1�!�ሮ,���k=�.D��U�v�E��Ң���g��d�O�9�tǳ�v����k��t����S^T^^4Q�����>@��SC�r��G����ф�+n�$Ђ���-,&��"Wk��@�|aK�������+�X��.V�y-�>�)�6dA�g�qE��&>M�ߣ��#p�{vy�.`�4�t�7���.��E��L��z�E��x�H�e��!B�ܩ{nET��Ҋ�K�����:H�NV$4vu���'�	��7S2��I7�"��LX��v7ſff��{�	;���{�]��>����._`U�U�D�8`xr�t�ruy�j��aD{�R�ۤO/��������G�V0��5��Gj�����f���՛1�Y�A�Ԝ�4�9��c�x�6�Ѽ��	��jg&�?�!f7�����?	d�E�Ȫ~U!���r�J2kur���3���]+��	��T�h���3��=�x�׏LUK%�:P�?����+�7�N������/�v��1YZ����1M�(�[K��Ɖ�����aD���2`ǣ�W�2����ط'5̬�2�}�T�aH���@8b��X���X��kD��Y/蕇���8�}�,��HzpY
�~�nd�[4�Y'�eQ���[������,��L񋾤-�o8=��Q��^�8� �BmZ�R7,���s��T���*�=�f�Hρ���$K��<����������}���W
ZY4P���AG�f�'�v;���S�5H�8+n�_O'ͻyJ��o��a��t6{O��bQ�qޘ�>�A�t�Zn�G�bq�4X�����������|���iU���f�nԅ,��k���ژ���x}x _��zP�f�7:1&����o�Ņ��d��U����к��N 2���A�❛�9� �8e�|���#�T�f$�D�޲e%�{z��w�aQ���
��Ї��j"����/�=go�]Dx��>�X�H`ٹY�3;S��%�Qͺ5�9�ƅ��-�L����@¯J�.��"����y���A�KY8u��]A�у��T �̽�o���S�����7��{��_Pl
�1"��I�Sk�������r��m�gh=[Q�?��,����8g*`�6���8��qi�紱l�f�mi�}�>}v"D(�Ec!"�UM��,mя?��.�� F������f�z�dz�<{{�,��G�R�G��W��]��h�8��#m�'u5���c	b��ޖ�<�� W���T!%�s�T@�k��_�)�"�>4���<��"�` �F��f����|՝��)�~��y��
�,;�脦c��p<e�K����;z���<�T=�2j�����fu0Q���s����=+�}Ԏ3�+�YÁ�\�0Wj(�!]\�C�`�p�����`�ݞ��9�9g��J�O�֕�N<����:Z��4Q�=�š����u��5���+M���P�����@`�V+��T}#��I) 6-V�!��(Yx;��5p�ԙ�{�X����ԟN�l| ��Jte�%����L���/�Va^�;qO�������DV�������9� bW�UGz��"Vp�.wz���#�V|M����T��:�\ݯ��=�����8J~Y�ؾmN�`v+����?��������^6J$��'�M�kGA�#Xt�-�y,N��8��2	�y����\�֐���m�h�qy��͍�t�O`eg�p��O@�]�S�:-�������;��%�b�!,�v�c0CG�XT��(�A�?~�:S��w����n�g=�]�!�����UK"i���ڗ����0�O<�$|�yb�v�b�z�D�5����ϱ�~ m=E0S|�l:x�N�|y)�L�,XS�X{��j[����1�y���%z�)+r����ce4ooP�T���^ǰ�tj��f�_�V�^YϜjUh��P��u����G;:��x�xm|a��^oNT���.����fj�LLM�B�=,����|j~�w�ڼ �L3'����{N���zlP$�kѓ싇A|��f�����ReMC��T�'Z�4��]������J��m6�Q�2̖���_�t���j��:�3�Qӳ�;�jRO}�V�����L�Bk9��߁0W��t{���$'�Ǿ�nJ;޹.�{�VQ��Z�H{��2;���F�����YN+Z*����Z�����H�� �+�A���k��Ó��p��&~l�aS(T�>�
����iҴ�ѡ��ݢ�"kӼ�׾��BL�rST,���Km�X���!��x�Gi���n;�0R�J�ކd�3�bZ���mJ"�◖�?1y�-h%,��)/֣(�t�`l�<�3����0��Ю(�>���mas/0���,P}�m��ۧv�8:d��ޮ��)�"�ߚ�{5��N{1��0�m`>Fx���D��%w9����?��kYE>�}�ͷ��Q�e?i/�e�@a�*�<��m����H/2���2aM�}�KaȨ�T�~�[nQ���Hs��}��ah]ڙ�N�O�"���7�/��]��0��&~�%$It�q��B>6=�#ڲ�n��8=�}��ʐ[y���֑A-y	�VcY��-�ۦ�C������t�)���Yˁi�
;X�n�,N�zaȠQ��d��¸^>]�_��o��K�'y�o�ʇ��W�E停,Wǚ&�Ԣ�
MH��p:�����]�y��;A=d�*8�I`��}��*%�i�2 q��PА�Ѧ�99N��j����|��S4Z?"��6{L+(��: s׹�*}*�`�fI�J �7De�J�;�#�Ǿ'%�b,�Y�RZ)<����k���4(_��f~��nb\/��f�0��gml��!H5.[OFE����%���H��MƭH�Ȇ��i&�}�z�X*�\*��\aHY��"���N�����\�g��J#��Lg�ʏ$�}�#���c��R'�6Ս�8�W��,Z��+�P&{/�[Xeco�5�[�RoR��4x�U��S� ��������?��b�u�If|��M�؎�4=� �J��������!���.,��ϛB��L�^3n!��0]-��ew�gP\�{������+T�g,��A�\tűa@6|?�1���+��ٸ��a��WBZ��]�����g`>̃��C�;���Z���+o���T�V\ƶA�E8���/�����m]*A?�	`�ҡP2^x_`�ó{�����3�d���o�OfpS�h���C)M�A��2�v�����1��?���e�h�I�ٔᬅ�)#jP'�"6�h"��xͤ��|���kI����Դ�A��Bꠦ�6_�4˧���~�&(V�>�/D�:��h�TW�bI��6���od&$�����5����1V�X��j�J'�}	/nm/�m*���ϫ�e���;Q��X��O��	j�F��[T�$�p' ��5
����o4;�^�'g��+y3�� $ƪ3�����O����e�`�+
Y� C�G˿1��`I)��}��\�C|��]DX�S�_]��i3����'�{Ip�3����N0Ѱ$#<�'����co	� 5��7䨠*IN��v�=�w�S�Y�h&����26~ ��]QZe�0 0I�}��]V���*��Y�,F�~^ۗ��d_�v���Z�Bw���G]X�Vd�[ b�L���{W_~�AP�����ti������Y~罣l��v�-�2��Ka�(�^_k�[!!�{�DK5���e�&(��C�,���붊�a����%�˚���Y7���Q��l�L�Rg �bǞtO�C! ����1*1M3�@�'���?L|�T;����nΔ�q
���2��Rv��ޤ9�;hmn�p%Ě}4�p��ʍ�>�l8������O�3K���UɾÔ�^�`db�gx���R$����Œ����j���w��$$%h ��#��3�ߝ���d�̄5,�51�J2�gN��| �׊��
�>{�G/=��4g%XR�[�r��$?/O3�M�'21=s�;��������<_��z�WT�A� Es�Y!|�	w&�U�J�L��3������K��6jt����Ň����Z�������'�2��8(�����~��b3j�!�.�	�����v��9\p���Ҁ���4֤�O`���0?��gC�5tY�{_$��T{�tH,������T(-��r�f��\��s�b��,��;�Pp��!�l��!ğt�TJ0M6�b������9 *�s3-h��6�����>i�	�p��:<�_���g	F麇�Ah�Qm����h��(mm�)��+by�c�Ȧ-�+МĆ��_錦kpU`�f����tav^���_Qe��EM�ڭ !q�B���6��@�:��, EW���|xNA��y+	���M�BzY��/b+�#�?so؏?����}@ ��8G�6��o�I��d��)�iӗ3b8Y���|��l1����$`���Wt��nc�t�����\��n��vB�j���ipq Hcw���g���b��|�J{��Μ����Y�����F���L�j�`��\4'�`�\�u���q)��B���y%Q�Ŧ�.�B�k�~s�4�""};�y�ڰ~=g�+W��f�t	�mxM<V2
����QD�<��S�LXk9�PrdՔ�w�q7eҌ#�=�� �x[L�_�+Xn�2�����h��c�x-��֨�$@3ɐ�)ˤ�k�ꝓ5�\��I$���������`�H2�g@����3�(􄋙�uً�`���v��X�z�r���ܼ��8������5Ŝ��x�� O-�(f���P������z���9]�Hx(�g9Ya5�Ϭ�%��3����Ȟ�0LĤ������)�>sD�m�.��b�3T��:V(���	��C�K��K- �BQ�f��G �f�e �w����%��݄&���K��|E�񱳫��[ìA���Y	�r:��E���Px4��$��[�L)�5�Gs�<��>o�j ٲOݫ��[�|��*~X ����d&���1�Q0G ���xe��֍�W�Qv� M�*̗/�`�R�V��7��!tў稾ШF+�s���%�N�2����(�N�p�p�� �r������h%��w�}�&m�����.�qfm�r}�����lRN�<�ֿ���!�PmaC����B���d�C�aU����ܡ�Ά��r�9����SX)����R	�<{�w0���q�˟W���ݴ�3��LBTM��~.��eg<��=m[�Wk%��[���6ֶ>?MȘ-��0�r=p�	�|�, ��Y+I*΢D�h^����ˤP�x�.�$���j��r��M��;�����1R�N�e�F��a�='�}�m����&m�T��|ƛ�X��yv�x���Y�T����5�x��-�_�d����� -�ध)uP�{oiR��s�ON]���ޭ��'V>IX��5��Q�?�/bW+r���mf���|t�o��p",�(����$�4e Q��)�)����Y$��v^�^�r�蚖��x�f.�d��V&aGf8�A���Ŭ�CV�AK��z�JU�]�P�3���Hr흚(��������@�`f�Z����5j�v:C|x*��#� ˠ��z?�4ǭ��x�:�ъ¹�
M���S�@@2��������=O�@��|��
��D�Y��a�m��/6@����� �`2zp���:'9�)2۾BI�3�k�x��*���p�IN��ڍ蘜U|����`�Ȥm|�%:���@9���B�,&0j��nMZ�V+��-��aJu�����ܗ`����R�#0�I�� ^d�j~ JB�0q!�3·���⇅^`E�N��L��i|�JNz���=C �+O�U�P����� �jllZ��h��`�!������j,Oj��ll�,+{[�:�k�ӞD�,��&��G0�B����^fn���Hl��1j�HS�I��S�8.��k~�`q��GWzM)pvE(�����?�eL��VU�l�N��4��е�⒇��_>ܵ��;�,M�ʻޘ�-������+��gÊyp��!���)΁��P��^�ʉG�7u�,�\�M,	��v���VN`�?���=�;D�=�$���b�.�vu!�/Q�MA�����3ʚ�/�VП[�{�Ѓ��Su�vB�u�K�y�R7�d%f����!��0і�՚�!Ѩ{�[i�D��2<g�����i5ڼ�ɱ��:5�B�W���>�2[U�Xt&���fE�왛L�>���
�6F/ۜ��I���ѯB����P���o2@�-���2IL�����Ni�{�&���$Q"?��=���Z�z����2�+-TTq�5�'O�޹tsq4��)!�<���lԴ�v������io�b/��WQKp��Uy5b���E�H�PTA�u7s�""�(q��
�
�ā
�	a�+����!krHPR��@��MLp
-��d&��w ���/������w4�k�c��$��Ny3I�}�}��e��4IP�^PD���ʉ���v���,�&�4���_��������h�"�޺?[�gٶ�s����ga�z/�����׻�|��X���
">��a�Ѕ%\G$wV�; ��:�v�ap2�1�>m�eA��h�PjVb?���׃6j����e]���uW9�`�H	@��t������[�����JPs�����$N�f��{��W�e�DI.QE����3Ըc�^8�m��N��#tH�y�3^xph�]h]���Dr}hZ�*�%�������T`ǝ	h�󻪇����<]5��p17�6����HW<"����YT���p�`L=����Nډ��6ho�?��\�C����	�h��j���&�:�����V=��3fH�����9��()$�B����5׭����H�L��=�.b�����X!
�gS�<�b��ԀSj/����tmg��ە��A�	�v�?L
�9v����XLK�[)��l��-���ѣ��VԑI�?�!���ih��^�/����h_�9n�9�[�A{���Íg�3�I+��]�ӕ��$=߻W-�����7��7-tz�AwaY����e;
���9;W��q�:\}�Z��L�f�R�{�F����\�M��?(+k��4���k�|PgE-�&�^q�-P�F�PZ�+���vb��T�c	nnZ6����d��l��ImUhݎ1��u�?:<^vmo�'{#�����s�w����I����}��Ŗ���2UȈ��':��:����Kp'�����Үt��m^�o�V�������a�ֽ�>�z�:�!�
�:%��HF�����C�����M� �6ū�j��N,��R�;�zHߟ���[Zѹ�NxQ?3V����;�����a3K�[�Ҋ �+i+Nu�Ŗ��[���p<��U ��������X�)�S��)L�{���HS~e��]�W�A�柨0���v1<b�#����,�������$3<9Z��°Ի$خ�@r_U����z�:.󱘸!8�(DaHt��B�U86��ȷ~��0ߩ4!�q%R���n����]�Q����RY�t`jk_M�SDLnJG���8��{O��<���n %���¬�����j딓������n�K^�:+c�����J��2��l�"h̭��E+��.Oq�ʟ㑽3�����X�6AV�2�Pq��#d6��.u��aA
(H�|;)T�:���1�����N�ވ���~niO���R*2�戸|�Q��E�Q���гr�js�$j#^'�O��,й������ �r� Us&�o����x;}u9��mjU�3���iNt4��\U�{����H;4�eb
җ��R�$�|�����h~�Ei��m���iHw��z��P�cCp=��6;�|�ѵ�oY��~��=.��tKp�I�N��Q�Y7� �p�:2�MPP��Z>a������}|�^�L��)jMb���Q?D�R��`�m�a�C�he���~��X�ۓ�xͣ&�D���?*t�S��F����>�9$R0 �b���HϹW;��`����H�I~y�} c�I�Y�-�ٷ_y'�Z�������D��؋�$���vvO(�Z����2��$�ԆKˢ���P1[s��������������hp�kqɀ�Η?d>7�(��c�d�+f�w�&�d�Ġ���+r��J���.��km�5�#�ƍ\$�����#K�Y��7��@�V\�C����\�Ѵ����L�\#ɰ��<�ZL��2��S$�]��?6I=�����-������7'��~�(���"W���bHP3.h���9oi�f��<��9}�	Ւ:�ꍳq���(�	��ՙ�i�����p�04�ao��!��YOo0������C�.w���Dc� ^kb:��_��l�T�E�nM	�s�O�[Q�X5N\�51O�5������qU�AE�M!�ڒ��i��b4L��<�)3�Ԧ��4��}��X���g}p�Mx�w'��V��V!����,]�-�\7^���3�	hDO�K����D�Dgn��(�7{�F�}X�pS�}W��n�? `;��I��0�?�'�8��D��7b^�����Mo���{JB������Cހ"Qe��̑d�,��ƎUF�H����w������n�$U��g�E,��;�{����  S���ؐ��Y*�K���=Z���ϩx���+��G�"Y�GN����TvF��S֍��m����d�-qu
s��^o��'�l�B�������Jj�jʌ�C�,��i�'Z�yJ�H�p����=��m���^�T]�	M���U���ί�q�����
#������a��P�<�]��ͦ���>z�S�[������ᑂ�.���
�"�}�g� Xj�?�#8 rP�y��_?�@M���M2�2D���2�~N{��W牁%D�b��ًp�FfK\:����x�Dó�:�¥�k!ѯ���܋���R�����W}l���m{���\c;�H�'��*��ڟ�R?�����3J��Ċ��'Ơ�X�66��_q
�}K+3g0�=
V�q���m4��׫Tt���ې���/�ڨ|uoOF��x����f;�������w�
����e��sb��_��!>�>���dij�Ʈ�ȁ��a����e�F� g���9��vy�޴�Em3���(S#ǚ�=��9����6�7� �̈́���a#t��g´���������_ˉ��!L��r:g�,	ԕ�<9��s����r��*��~2���J�[Ś�0{^+t!�� `���"�`F���>u��&�K�r��=�D#2�e���Epƙ�7��H�~W����+/����#3..�	 ��Z	J���('SS���}&�E��@�"�V�X�w1.B��Qʵ�`�,n�6d��R,|����~fȄNa�=xa��D;2�8f��4̮�ׇ�h�%�=0d�%&G)�Z�_�w��e��z� �]�x�l��%�"D��5P��Er0�J]ee�NQg�(�_����;;XE��x���t�#1@11�(yƸ�4��@k�P���;���z��c���/��B�^J	���Q��@�9axI�>5օ cV�;�l���0�!�'�@ӈ{�P��d��[��^��J7��1��?l��=܁|b%	_�ɀ����Ż>�"D5�GÛ E�8o��T�v ���FS�֗`�$����$.�\R)����i�O�rbRiM��cP?�K,�m*�{������C暫��t�e�����0��Ʈ�I�(�oJ�sǇ7y��͝��%�D9��:���h+��Mos��9��k�i��+��,MZЇ���� �u�a��䲇�Q��x�,���,�6�+Y�֖��T���U1��	.v{�*�H�����s�r��Y�w7�=0�L��F�HU�GaN	\����k��rTp�ԇ����������h�j〪�z'�N���R�/����+�ub��iEn��{�n� (�߲+{���A���e|���m��{��j���a��م�A�?`�mG��w$�Z�nW_�ֺz�������cZ�t�_5ɡtL�@�؆���_|ML]���I��:Zƪ�|G#��]&a���X��	���� DT�������{�<����
����>U�a��>�
���2��:]��<t��~�p#j�񕱘×"��	Z�˗�;ʘg� �Ը��#ļufE�����j5$4�cX���ч��'C
Bǔk:X���|R*)/x���� $����-#��+�@�M�/}��!��
�U�Z5�uS	���]$��9;vvO�X)Cì�Z�ڍ����baT��׼i�*_�Ui�k�J�iP��$���2Qa�u�[NĬ�e���Jcڦl*�( �4�\=[9�Sy�<�ϥA�8��zk�)���FX����C/��������cX��#��]�"N���O:_y�o������<���q���1��S>�'_i驓5����XbT��R$秊�^���=)���?'R���(Ɓ'.�W�D�#�S��eh��P�ST�W�r� <9��/g��'X �4�m���=��r_>7V=Y����D����L�l�����D�(�DJ�����Ѹ䏷1�	���x^JI�R)�+���8^��n��(.�v��P��(�Yu��w����׻ź��g�jV�$�8�VUr��<Z�Ƶ�I3&��R��� v#:���"r	�i��$_	������Z��m�#߂����/��|\���=���S�&�l�
�;�q�&�K[CL�VmN�����Cϲ��g�U}J�ס��@u�/l�d��):�&�a��mwI�$jv��.	R���qϯg��eI헀 D0͝P��8�|E�����=��܆�U�z�5���w-N��%&������kV�\Ƽċ��\E�C�xf}�4I�aۜH9 1ܾa�S>q!)R�w,!�j�U�6�5�+wmNX�^E�w.ƏP��x]8\&��ܢ�Dj�̐ TZt}@��'�����z��
}���B�V�ѭ�l��x�Ɗ(���a\�$P!X�L��Qj�7s�%L��<���ohH.u��1�,�	� �S:�����g�����s��v�tP2h:>��=�c5,�@��31�9�rDY��){�[̱58��✆�	+�C�lc�7�9l����ےh��� �X�3�m�
�Z�9?|x�N��K�6����]T9�e��6��<_���%#��J(͔����dDK~�z�����c�U(����'�k�*.|%bf�F�{Re�HG=~���ͬ`�ܠ�k?���M��̝0�3������	#������ޤ���dFR_���b=�P�/'�%���.���yd�$�'���BXB�$�R�S֩lc��Aז�B%��$����H%5��p�L����7'c�L:�ڣ�럦b->9��g�0���z��G�M`��2��^C!�G�Iߑ!#��=�������o�E� 3򕲹�!K���d/���s�?�O�l��vWK69�ҙ���;��y�9�JO�Vl�F��u���p��Wֵ�9��0OB�R
�sBQ�0*oJ|f��~�Q-�(�Kfl�B-#���{3����4|�\:�+O���k3ߴ'��Ef�f�w �� �,�2_X@��"�=/ǀ���ߞ�eouR����۟b*ͽ[hS�Z
�I����������_��H)��Z"�z�%���ܬ�"�ɤ
�S^e���t�>�M�>}�ڈ�zm�	����KO�y��#��٤a �k���V�囪��$}R��)�5`��[���}Ӏ2T+��>�}@i_L
�3z,��&��hjO� ��k@��7Jˢؕ�ZވIj�j�"i�z$������`3'�{�<�dj��Mt����Ġiǵ�� ��'�5+� ;Dd��`7��ͰH<s��&@���)�/��_6��00�]��l�b�=x�,פ���a�訡���Y1�脂tv���ҙcZ��vߦ�)��r#'�i�Z��-�c1�WK���
��v���ӷ(H���S��|M�9�*U�@!���=g,�K&{�V����&|�o"�MA�=�eyp���E�Q�]���}�i��ǒ `��k��讜I��⇟�r0�3"�?��)h�Q^U<zy���hX@���F����C�_9+�DY�@1��p�D����C۹/�%D%�EJ$2��@S���p��,J���`���d�%.�����k�[����9�&��[se#?':�(>�2���7@ײ���w�հ�V��n�b.�w�����1�E~y���6��n�.�!r#�ޜț.��6��1O׻�$5�Q��~ȣ�m����Z/�S4#�|���|���2h��(y���x,��!�m(��<U�Q�Op'�k���c>c���~Y$ 2�t��V�s����!.b%��e��6�������wV�G.vk&����-o��;��~��P�T�s�Ђ)����X�Ȇ2��؋��*{����m4�ꟶc��ʿA�N�\V�|���<LE�A�V�ЍJ�����-��&�{�0��I�8�<�q>�i5 I�k�'2Mҋ�ac�RP���Y4�5^��c�y�v�͈�3�ͬ��S[�tFl�w��0�/���G{'l��t[T��ٰ�K;��Dg���q�[����
	S#�gC�MZ���n���y\A�G*�E��dv�W��Ό9� 1�&ud�8G��/��ɛq���j�؎��
"���y���Mr�Ӷ�;/�I����i_�N]��5@,��rI�T�?- A~J�l���J1�s��N�ug��.��"��G �n�0)*�=q�7�>8HN@j*h�/L�&[4T�z�#Ӫ���a�aI1�'���]ca�G[8�oہ�b'!x H��4x���6l��0��g���!S���z�B	v��M��5.��ې����I��`���`��7PMc��-fg�_٬� G���D�s�#��C��D�Y�u�c�_xd��vb�c����JZ��=��] 1�]�V�XF����8�C[�������Ϟ��"��.(D} ߼��Nέ�ޜ���0{;���5G�ۉ͹�}�����h�pH�j0 o�q5M�Z��F�:�6ߖv"�.2� v��V���vǞ%ngM��I���wc�4r!*��U&�ӫ?���Č+�q�zF��sQ�:����G�ئ^I	OLN/�M-�%��g�N
Ug8�K��!b���-�cxX�E��+we;�����	�1����H3�>\><{�e��s�]; :��P�	�� �B\$`G�;�"R	?�AO�O�ی���ཱིNU]����`3�� ��}�"��)W�=����!�;���M�mVʱ��DB�PƬ����F�\K�ԣ߫���f5����R����ā,1\E���#� �Y�k�y���Os�Ñg�[.Y�n��_�`ܡ.��4Yd6"�tɽ���~��
2��e֎ڠ�hn%j>�o_�=
��Ҏ��:[��oh�N�����G�krU�fk�~���H;�YI
��4�������� @�G�Q�(cA���/�M����w���l�5jYD����:C��ʑ!���j�R���"s�z	��_�E��3�Y��"L0'*��\��b�b���F1ά�_Y�w7:sNr�������v��ܣ�5�ti��:&c�ۦۭ�_t;�x-�����fdᮕ�?ۙl���B�z��Y��~ߔ���h�'>�&�� �ȞSS���T:�_ۂv���#���U_Ňxfdb�f .��y��p�tC�}��bz�*.z�pUXwڠ����WJ����zF��;0`�DC����S��g>.�ٖ�ͱI�[Y[kp����Z�cn����]���2����f����7G���>�Գ�F���OYyR�G���"ݵ9g���F�7�: `��yF���*���`E'����K�+��p����eߺ�����Ѻ�>���WU[��_��C G��\����g0y'P����的%AG����H�� =u�9?��v6�3H
�+�=�Y��؍]_�Y�D�JI'ҩm�%A�"C����Ə.xx��Lh�̌�B�`��8�F�,>�!�Kd��-}�%�
�vj1u.�f�Jұ{�ni�w��h�]Ӱ�~�0}6&o�[Z-�#���o��ݭ�q<����=����ZEyŰgϖ;DJ�S��'2�:���������5/���3'��|���:�n���zB`�¯kj�7����*���P��΀�GN�&R!��=
�I��b�绷U8�@90Z�|[~�j��(�lIo:�f,h�s�q��W��k�~��C^.%_�|�@Z8#4ڴK���'{��Z��*�Q���Pm����G�yKi4�K`�+�*Qh���.bq�@=�	�tS���AN�����d=�P�Ɓ��a<;2���
�nۚ��w�<UtJ P��\���䡠@g�k��ﰻ�Q&�:�H��Иi��h����]�!C�M8���S�p�"��d ���Q�0���G��-ۺ[}�<(�4-<����r60j�*�)����bJg����)w�����^]���j��P:�v��ThGQ)k��(�Ge绬UCP���Ԋ��U�Ȼۛ1Z�a�+�6b4���
�2�b|��HT�Ĳ���8�T�GfE���g2�0���K�����ʃ��0��x�R����y3�G��q-��]�=k��f�`�Q/9f�qq#+$r�:�Js`9�c��E�{����C�4ٺ@�s�xW��S��Q��
��N����4˷Ax5J�	|�\z:�u��p?��>�n�o�VqIj��kJ�l��LQ`�Q$�dTq��H��!v[�p'��7�����׀��,�SW5��}f7��R�KS���41�Z�G��u����_��I��C���V�`�;��&����o���ÇS�h��Lhq 1F.Fg�qo������m�vr��˸g�&��?nru���c�IV�4���2��t:@w~q&q��_�Bt�V�����El������Lwlϐ��2x�fΣ�1��F-�P�?������J����8P�&�t+s�jg�L `�+RVǯ�6@��	�}���e�W-�qd��AJH��#o�����h�"_F[�<O� ݴ�Nf/k�"3�$���.K&�p����zU��"����8�������b��� R&�;��iԠ�Ym��8t �����; ]D[7k���5"���\�ͤ�wa��7Mv7��t	AEB���dB�U9Y-���$��0l��S�i�D8 ������`%����!B,X�^t�O��Z���sk��uN��l����,�;KA��.�;-7YB�3�'ߥv#�l��j��V#k�Eڲ�[��>�Ⱦyy7\K��9n1.��Q-��*��>�T	LԼy����!���;X�l��`��*�����ٚ�r��HO�>�"�&��)B�]����G�
�A�� �M�{`%y֦�@ʭ�����h��h�Apq�l~��v���J������D���X��Glv�Y���*uw��F+�<�a�è���ӓ�By�_J�cG�I�c&�x�Mƾ^�=�s�3_��7��i/r�¼aKcs��/W��	���x+�A�l�����_�ɸ �N�/���E#�-V\x3�+� v��4�Ù���]���^�lc�`7_69'�^�w�X=�,p}*���^�7���y���I&�����<{y�/�l�*���&��c͹K<^>�f�?2�ZZ�%,��fO��M���V���g%o�s�!�]o���]����y����顗�ה������L���"-�'4�7��it\�H��T�\�����rah�P�����\#�pD
�DI������S���8�n|+�%��'H������H��{���;��A�+A.�hU��0���E��;��*Eb� ?�+�#;տ[�Y#�q� <c�4B�\z���,�P� ��3�n���(��kv�x�w�b�v�a8�Ǘ{����tB�g�`�K�<`��+���~���=�]�~7���/�4��k�c������d	lP`���YS����O�v��z��ٚ�-I����.r:�k���/�O{]�<�����E\�ǜ�*�8e,��gLoϪ�x��?�|,w-���[��{�Ԭ�x�J�ꗦI;�x+)�'_9�n�x ��H];0#�L-���BEX`���3�;��_����nw�-��&���V�[��IMJZq��l-��R;���>nX'.�T��E�����A�B���
6�
�L@̫dI)
���D���Ѝ��z�M���c+�3�/"�|���^b�K��� �<y�TFK�b�X�Pm`� ���_l�n�+��#S
]�%��i�klh�=&�/uº�G.�Im>2]��(���k�]����A3�䀹x+�TS�����?,�E ����&��9�+�¦�+���=P�	���m�v��kMQs����2��w����\S�!U_dZ_3$L+�/��`��mY��"w�M|U�*(�zI��@����,��(E��E9
��\3'>���h�]��r%�g����II���i|گ��v^B�=�>x���?�k7r���&��.��f|Ev5q>��b*�v��w��T}��S������wJ`v,�J �#Jگ�^�^��.���\H���a�����g�]����C�%'2�
i�Qt-7KG��~n|��
�w��͕d�. ��ea�K��
i��:S%゛���"�C{�Փ2-+$�nls]G��
�,2������i�f�ruc�j`5]wY�;��Z��K�׵25V���c�κϢ�d�R��#X���@�O)܋6&������:&(}�l�@�D�>��[-Ao�u�8��PM�5L�'�w����hOG�Y1�Aq�Ҽ�����6-�y�аf�3M��u%tW˶�#����uNW؁���_+�W�Uq�)��;����]�ǫ��l�dU)Z�����.V� ����1��B�m�z�#�-I����.n�@F�r���y
�MF�(l~Ǉʡa�˂ׄ�Y�^zxt�f�-%��RЖpJ�5�bǇnr�SK+�W�g��,�O5�E-�h<
���h(��qlOTn�[�=�'u4+wx\�拾 F)m7�^�ʌ`���&��ࣗ������8����mS<̱������$������$Wkֺf�����r&c� ��>:���Ȇr�R�K��nZgp��_��gs�o�;?��Q~�\x�Bs�l�"��O~ 5x~���0��	n����K'���p��#���&#��A�EMiǸ�Q���M��_�B�T���W�f*�;��2w�/�I�)��\וs\V�*lo`23BD4��L���Cvw��!=�T5��p�������9Fg��X����d!�����8�C���y���%�a�fi�%�κ��]P���g^&t�:kFe�;�e�N\\�~���2|R;�N5��j����՞��.p�ti� ^��]W��|Hm���<�Z)�rpXlS����4X(��ч�b��84|�ݯ����!��:&��bw����v��X9^�߽;1�H �sB>Dhf�d���1o�S�I��aɫ�6�����CN[N�����&�� k2��=��Q2���y�'X}h�rIs;˳���0��00��a�k8�c&�5?i����Jq`0YBJ�4Gh��W%W�0�E'X�ݧ�Y�
�X�H�$?�0xy>2k3�F���jd���[�(}��ZmKa���\�X$�d�{����g�75g�IK{jl�h)aU�.��R�G� X�w_ޅ�;�рJ�%3�~�Y���x�N�৵���/g���UѾ��Ճ�\T]�}����| λ����m���p���('�7�?�w&�`���;RsAz((��T�緡���~��w!s����]r����z�4g2A2�2j!�Rdq��[�ֿ")�t�!G���EWTPZ�����ӓvM"�[+_�8�(���zo��o�����Uԏb% �>��ׯ�M��W��W3��陮��m��*�buB�QY��1��A
�+���y_SQ�v���w�]]��X����4g�1���RL�y�c�V�&��s�?4�*)��F��
��xhr��h%xzOn�i˪�(�	8��|�B�}�%sG�E#�Q\킧�Z9��n�J��ڵAe"IS����訡OEG���������r*n���E�Dy4{ı(EJu��~T�)0��
^v�OѲ��ZЈ2E �Bv�<�"u'�`������=�i����z�1�i�y���c���b��ƀ�?��������qQ�����J��\n�q4� Ōf9��J����UA��Cf N����0�zJ q_��ROP���I�?� �h�lV��H27�G��)�G	��ÔB��Y���4�,������-_����M�m�*�I]8�7��nf9��cF�-��*��3�<��-כ�웩R��K�#��hw4�1��d��ή��Nz~�¾ӊ9B���1*�`���,Ъ���/���_y�}vf�����';���B�M�ު��l�6�L���p��>��h:
=gr�+�=�Zئ��S��s���6�����>����,=Hj�	b�� %����s�n��q�'�"�Ho��V�Bf�z��J���\3{g��,�N��X���u��ru��\HT�w=(#�C����<�(�]�qK��A�`?6���s��rz�]�����{�$n��Ȋ)W�g�PC�-�+�Z�F��p0|���E��p���j���ۦ�g��D�S����^�ט�6h�K?�X��'2�bj��ܹ}�W��j���}	��Z�9�<PQ"(�n���3��T4�'@�Y���eg�=��3��62�I�&�.Q���qfk'���#��P=����T,�X�W�x�����"[��r�%��\���1|]���"�O�L�!��2��Q&�S�M��y\�Q!;��1�����3P�GC���g��������w8��9��B�~?�����6��]��3� |��[ ����MH��ʩ���N+���xzM�����c(v�&�U󐆷
�͘?	۾C��4-�O����X1���]���]�G�����<�:��a4��N�'If?i�7K�L%-�!8�n���-8���n]]d������O�3�Qy"�я��/���P�}��+r�_Ϣ�]�rMM�,�V��0�EK�?��j��j<�q�bƔr��l�%� �����$F-dy/<m")?_xn�����l�|9��={��6�q��e��ח:x�g�f]�mT��um�C9��#r�̭d��\E\6x:!ڕ��L����p�<�e��=��Ȕ����w���m�|�6��7ף�F��[:��ړ�Ob${���J�z�&�K��>��ڄ_�����m����.�B��L�9�1�䳂��3�Ƴi�[�^�0A~�-�����3������s�y�Hw��n���������^�v�x�-1Lj��?�@sK�s=O���y��8sB�����/�� Y��[3���8�
��;���#�8&UJ	�� %�U3W�0L�%�(�'��ޯv����q��\L�J�:�XQxJdG���Y5I���1wJ�'@a�u�K��,�	e�$Vz�<T���[e3r���pϰؤ�5]R�5�J%�|!^���f�{� �N�x�N�ĳ;%օ��M�2�fNaS����sщ9�@'���U�z�T.Y�P!�b���<#w5��[0~�?�5�#�k����|W��?E�����Zk�@�˶RHWs�JX��&V1��{_(�N&�(�M��M�3�
��&wc!����֧9uX�M�Sgnu�8起(k�OQ�� ��j�����"k/s�gv�S'�Z����q�Q�	��$�A#�	)�<cs��}D���91�\��d?G�.�Ks��{��q����h���'{�}��є�Kt� #���:�M�����V/yF�&ڱx#e]z���C
���6ݺ���h�i)={"�Di����?𸩺"��w�}�GR�����|S����%��(ٶ�j�s ���%E�B�iɉ(e�Q7��B����{�ť��Pg����t 	s��<{�g<�N>���I����":�V��Mړ�4�-��Ȣ�g$�V�Ywׄ�|���z0�66�a���~s��<8�ix��T�Oh;����%�U�~��']�����+�H���Xp�n]�x��Xg�e=��*-Zw�ZDl�������3%K��^��=�����ɋA3r��x�!��Y�V�:���LK`PI�(�Ƌ�=�:���~��ġ�3���ɚB��9���IQ6�]���f���KE`+/1���D�`/��8�]���Q%��*9�1h������ѐ�l��C��a��>�[�1��E�R� 5&���˺s�HrHV[HQڹ��QC�y\�գ��US�����9�OK4��Up�^C�"J\�u�L�!�2�v�g�$"��l*��s�ڛ��1���4��;��Y2T�A�_�{l�� ��eC�.�`߉��ʷ(�	e�8CGv���|��+"0'*�Y���|M��T=�k�+�����BB4�7"���p�	�-�`�O�R�j��M��h��,�{�T,�̳��1�`��M�^OI�Y�TTYS�p�cÙ6_�[��
� ;�	L r�>ҵ���-O�P�ͿuY��!ַe�����������t:��7��o	皞�g}Iq�&X��Q�R�[��p�����D���4�[f�z�d,�B�n|acF�#�����:C[(�Ar��d�:���$��7S���/�t�o��H:�����Z���^��Ou#������`��:�,{qiN�X.��I����#yuu��M%ȋ�y}�oiYm�F��fo`np��uߢ�\�v�z���A)�bZ����3ZJ �Ѣ-�u7��A�y̵�&��)�a�p�X�J}B���*��W���V���� �Z<��M:��z�[����C�=��������8�w���4��	C�s��T�u�@VÙ�I-Zh�01$�˫b�6���KC�Z��D���$�����ԔN�Z�G_�a����RYDg(ί��ũ�?fT!�C����Ty[����K�h5��˞�����m�;_o����p�0��,��\Qq�����<ɯmkz�1��u�H�>�!a��hI��p�6c�u�s�ڝ�����n����hR��rk��f����X�p �4�,�s��<`�(��q; ytB�"�Γ��|Cg��:A��n���P�]���b��'�z*@
h�2[���	o=�n�U0SC��+_��L�
��S�EKED*aZ�z��֖H�\���2b=����`	�|W1;�[ 1����m)��8����k�@LѧIҿ��u��/6o�R�kS�o�xW�5�_�жq���i#���_ʐw3Ң�D�6��YBau�	R��P�B��k�^��S���^|ƀ������'�BS�_[�=]}���|���^��}��0Ϛ+eW:da����o�ύ�lٲ��4#�a-�맫��Q�-#��r�%
7^-M`���7fhK^??Y�-2�i���C�*����@���J¹��m�=�A3��s����W1C��s���D�Z�j5�A�A��󙾩!�l�/�����K��h�R���>�)�z��4T�4C�P��(��D���q��G�����L�60�qf�S<K�kx	�X>QY����>ƻ�k[!�C�I�J�5Y��nE;��A�hˁ�&�.KU�U�'�0�sjD,�Y�o�!&Y^�YjU�����W�Y�r.l���~�����ǉy>�'���D��`��\Nm��|S 7��)9a�dβe�kۈ�F��k_Q0�l|�����Y�ڥ1o}����X8gع�ŋ���|Z+.^��o ugB!�_�q�?������r�z{v��5�*����4�ҫ��~N�y,%p!����}@�J�3�� f[H:	��4D���*���2�T���~�v��[H��Y���f�o��4�)� �U����]Q��=ӊ��
�a����:���Q/�^��R�����J�W�Fq�l�)���M���Yg�hVdW����N�x�]��%��j��I{˘Pr'V3kls�g�@ƻ����Jy�G�?��q�ݗ�_`;�32H׏A�'$�T���p
;�tM���pH��-C��}��-��MC�����u���a��rA��1���E�b+�3E$�~a�W��x�qm��
��/T��"�A>R$���p}��c�|�lL�/�z��N@l�vɂ?b�l�f��
�T'����;$�K�U�*�:W�ng���#.u�ر���	{;X9I��d�<��$�{[g�JY2���Ð`��7語4RfQ��\�������EH9c����Pi�����/s_�#���	5_�W�ƻS�6h	=�3�#�I���
���j��yewAC��,t�ܑ�E'	$}s�����#�l��P�ڨ�8&j>Ќ��P��L���K!S�u��=��~ ��ۑ����<T�Q2�%�z�gC������7>�e�$�w�Ղ�!`;6^੼��t�L'y{����QaS+\S�O}[��}H=A���P�-c:�d� 7�j$_W&4�2e)�V]�ո����.�a�C+⿲Ҳ������N��j�M �����2�@�Mn͋�[�8Jt��������@]���t��F�.%��C޴x+�K,�ıH/X%T8�ىN��V8�j2����CGbܣ{QPw�A�`�Vd��u��U6�����C���kL�mH��l�,{Ly/�5[�h�`@3P]�� �)X�Z�J�_�E:�R�_'��22iB~<5{�+�i-j{j|'�遢�x����Ou˾��Y"�>��N���~�*�Q�&�e�}��^���!L�$�-��S]���8v�I���mw*wUT�Rʚ��-en_z�|5ȿ`]�܏6kQ\�.��Y �#�������&�i�|_\xX�u��	�|�	-L�C��*�����)�ZO�@Vש�n�Ѣ����^���N�T�.
���,**���}�(h�w)���N�a��"Q����0��w$M��c�&J��@զF�햍�˄�c��js�л�b�7�������N��,���8[��᝘�4n3^�3�5����D��t����3��������ɉK����MH��'��v��w� ɿ�P�q��(gN��i�35B��l��͍��d����^����Ψ��>��^���
�타����n��ߥ�8몱�^:ֺ���K�B�'�I5��\| �jhf+�V@����"�ϊ�T�0�j�f���7���yq0K9�&����#j��l�=.��>7�١q����P���|V\a�~rE�pO6�j�]k����F^5��H�ϋ��\���q����?��&�B�>�"O4��.����d=kB��^8�䣱�p?Q9����5+��g�'辑p2�=L�b*�)'�C 跿����p���y�O�LS��i�A��9��Eޮ����n=ɡ���L�&�1��R��2z��*��۠�i�]���i��(�����	��9�4��)=4˫�f�/?�e ��5�"�*��	mz�#%:0���� =s��,�prܱ�	t��/���g��t��HE��a���B���r�oNp%עOd�c��m�e���V	�HI����~@�b�y����:�<F[�7 ~L���(v�"��0��a"�uO8/	qYh��O��Z�dt��<���q��>�����>,���_�R{���Y��Uf���?f��*lc�
X[�2������g<��7�6'���� ѥMX�	�x{+��,
�L�e�EɹZ-�2���n���2&�K���Y����I
���b)��՟�Π_t���EM}�ܧ�4X�7�%)&,䘴{�D���9��$R�r�B�ȨJ��X��4y��J�'*�M�&�kE�jJB|�2i�D�=_ۮL�#ڲA���Y_>���1P��������ۻn���������6ٌ	���`�b��C.vE�Hm���:/?���t�m��#$/�ۥ�П��jD����v+O�d�f+�V���G�� ~>��æ4�m���/V�i^�(���jp����	\Y0�x'�͠K��e��Z�m5��W��L ��'�d!��(���]�r�	�q�Ǌ&���×*�X�����E=鏍gq�-�xX�F͓|k�7����]m,���*�c����0�}��(��<ȿe�Fq�@�@���~;�����x��A�|�ϐ4�� ��В�B]1���/1{ԧ��ѢV����x�b��	�U��[@�2[��O����~�
Vl\4�BTI���M&o�;����^�V��5N�w ^T�g�y;:d�2n�.�����?d�9{c�70(����֬.��n�<z�}ʦ�Q�2%���Fp�.C�.Ov;pGk��DI�U� �9�k��K�E�G{�!J�eD�f�{N�g��� z�x��K�b�z��D�cy/���8;qG�c�|�~Js(LW-�e��wdj݁��N��s���Ƽ�UҒ�v�%��{f�����{h-z�������&��3��u�<8�����d(� 
a�$S��_^��n�Ev�6��$߁�� hd��v�B*:;�����3q3ѿ1���JGF�t�k���K-�m�6E
����7������-�<��݅D� ��4��vq�_Zı=]��K��v�asg��[�N���tu�����6,�3C��>]M@�C=��0�鑘�&�c����Ea}y������fPweH���NN�\xd�����"A�e�;Ih� .�b�~	*�_I���GK���|��T�!�ٿo��6�._B�=�r�u���Xo���ή�qѪ�5�}���;=:��	��h�D��UL�-&r4�8���l�O�w�TC��vE>�A/}���:����a!��P`�*0�{�Z���ע#�顾W���LUp�ÕW��
Z�ʔ�	a�N�4�0� =��NN��a��C�Җuà�0J%Cb7'����|����Ok�D���9.-~�e��R[ҟ�Yc`7C�Z�'���n�;��n�Z��jf4�H�N�)	֛����Y�(^�~�]h۟q+�����`
�]�*#�$Q�� �{2���dg�.�A��`�/~��L��_��2�3��Nm�}��x�VBV�f8�0=�'[<)�s�U=���K�����o��23=��KO�q��n��fkd��j(�}
 �s��QScE�Ԓ���E(#����S~-�"v�K7�9�G�hu��]�#
��a��]ǒ �[�DϿ�	r�ʧsdV����N*sz{�6�a�Ar�<ҏ�_�vp||b�M�6Y�:w����O=o4M=�{��ʘ,�_��������KK�ظ�s� J#J��(��K����&)�S��l,p�M��d����8�h��~�����@�ݧx�s�*0�%�q�:8Ʉ��r��r3)VB���6W�i(?Ŵ᪻�w�m8^������EvF!ڶ��Ԙw�3�		E ��������9]�\C�� x�/�"����;$�.4_-�rt���+&qț܆�t��MB����7W��[���	0y�e���J�my.�j�w�r�[z�O��[9�@��R=���	T��~���v��韱��qVW��{Й��;A��#`�`����^�i�]�YDm��Xh�`���mikKӺF5��
��Z��:`����i�!�U�sU����R�r=�%�Y$ʢQ���f��a*�����:��Gm?Eb�u�{n��l\�$�C��x�H�E�bP�l�u�S"�Ot��T��"V#��:�����ް֔���Y}1���9��;*�w�F�F�}a�É��A�����<@�
�c���Sx��(g�l��6����R�݅�L��WH���kY*�E��� ݿ�������D"O�<��"�~������JU�#�j`&T������a�t�����֡��H�2k ����n7�����c�a��g�׉/�x{��?l��G���<�cC9���_+#.8?q5�UMV��D#.����TЛ����U��/"~�}�}5�. �m�f����A��՛Q �ݲ|�s|��#��l,�+��b�ȓ�{
�� ��}����&�hn�Wc���XbW��y��TsfV2x��܊����ѹ��β�$>\\R����Zm�3haw�����y�G�����5.�h7�b�8�v>A�����B>�t֪�T���\)��O��\�Q󳐁��\�ዊc'e�m��d�H2�8�ݛ�dw��ԟ��Τ��.�矜�*���L�M�jL��(Ml;/3pq�,�́��:�/g�!��};fQ�L>�P� ��HqF�mD�����с�ð=��`fa�l���R%�z,�W��!�8ֵ}��|ɑƵ�dg�
2�j���WV��/$Z�ģ�4,/\���tѧ�l~�B܃�i*|�5��_cj�|Uv��Y�2� +��ߗ�&�3(�1�b}�����w�4,�?b�`�t$�O&.�c��G��8Y��6J~;e��3���S˥��pr�xg�}���/����*J`Bvl2�$��#6�]U*��o��RJzk/�N(6�31Z�=�D��|�(�ػI؃R'��j�qz��6���ׇ�ܫS\��}G��Cw8�xL��!�!P����j��������c�$�U���ҧd#=M���`*ā��!he|9iTFĻ��Uy��]�
�%d���Ar��CĢc�&l�r��[�>�Sd�kk�b+HF�AN5�]z�Û��[��K���R�Tl	�z��(��v�Fp-G8���5MM��1��E�N>��j�Y7�
nؘ�>J�`��i�����u�����������ӽ�(_��{,5��H�R�*@.\���j}���}N�Z�}b���iH��f9���p�����w�a^q'��5������]F�4B�z9kg�~�C�]�{TE3��&�h�7���tN��7/�cn-�de��>�/�.�Dn緰��rs����mR�$&v2�I
��fXa;������Y��1���Kт{��yg5��"[?z�Q:�Uo�l迿��|�2ՎZQ�U�A��c$��h��f����ԥ��t=���4e�iP|��:(�Q\�,	����B�GW7��)�F;�Z겾��Z|�g\[d�; �~�	��n�x e����M�ۤ�}E�ȳ6�fs,��x@�߫o[��'�li=��/����$�%�D��jk�Z�����b��Sz�z +����Į��9�o��N%�x>{���m�t5�
�H��`��CZރ!:����L�t��h�%6y)�)a�+R�vR��g�FT���A'r�+��B�`��_���v���D���O[����**.)�bP��[�;��B��Q�F�$_!�6K�L�KGLd�i����Ň�F*�Y0E�I���II���.�p*�ig�S��]���tD��G{+��^����5�)��gˮ�]h����c�M|1��O�ƛ_e�d�����
��y�h�B#|-J{E{fo$�5��W$�#֩�Zr�D�[I>����<Q�GP3T
S��*�1�;�MۿD�\�5Cl��[uW�@���a����)xӤ�;�7]k���r��A�	o�� -��r���?��nD�@����s���Ǜ���t���}��Oԇ�ɯ5~C_rS(O8�̍����܈�����1���!�����Y���؆�m4�%�����#�dn��7��Y)C������T�/�%��Z̮E6N/�О|�����_�ܽ˴���s3U�t�kW}�ty�ϟDxᣕ��)yk=\����J��U페7Ѵ�,����L�in��Ê�Z��qD��IF�V�"\��[_Ngȃ�7yJ0�Er����^���jc^l�����~	klw�����@�eI]�X�K��zS{.�v�[p,��K�9�۟n,�RS�_�g �ڄȐn��pr���q��R�uP�HÌ�	�[)VD]��6�V=���%����R+����E�00���ښ���t���dS��V�1�w]ra�����Q��'~6B�e�EB��#��~��S�L��/�vh#w��?!��h6���4��Dx�F����� <T�K��T>�i����x׼0а�b�}��7.}u�^S�ҫ�#O��wwO{��I��Go�g����BV�]M%r�_o*�c�97k�0b��Xa�0^��讟�.r2^n+J�KS~�����t4�Ѥ4,\! B������=���9)�ѼMu�Z�VU�RȪj$L�����q���`����ь&^m�#�`]tX�*?&U������l|��;�0��N�Q=5Ȣ㨜�;;��h�;k���5�$j�6�a��k<?Z�����2��)���ahG':Gċ�Y�0��s��kiZh\O���^��W�Z7��N�+��j��������Q�$�� ����
�TB�c�y�诫�=�[Dm�:���l�?i����km%��Έ�*�!��Su��N�؀��u$D�P�dq�@��,�..0�-��J ����V,���И�<��V.hJJ_r�uu�x��Vk)k�Mm-�Q�wZO?�M�e !���~�+��\�h�k1ɟ��ڹ�{4ۋ�B�J�����pA��wsj�s/��A@�/�ZE��d���fR+��5t�1Э�G��S�Wj�
�~��	��)|���n�9a�8�F07 ]�����D�
��ݷ�g�#�ә�����M��Aԛm����BG�v��+ ��&70�f�)�����J9��f-g@�VC���4aZ����������9�|�LػuQ$�y0=�C;�U���3�羚Z7C�1�=������O�t8lg]Bk�|?:��5M�AĬ+��%�g�6b�'����ZCPY�.[�>�w�������]������2\!KN�GS��n����m����5Wl�bEєq3�S~2e��i`�� �� 6�CF���7���$Q�*���*2�����~�i�La5���i��'�uq/�+!D 7�0��U���P,g���HAh+	kA��5��/P�5=��4[�j���>����I�}��i�b-���Le�!���֊��7��y�/`�7��~�@�!����F2�(B`��+�зe�J��",-K��#�E]��b�ֽ��*Jk�鸏��
>����I�ٸ���KK���;�~w�������E�=�g��/k�p o�U�9>n�����QM����Eе�����1z7�C¡b�?8����r`�����E�$�CA.w�	�q+_� �[��SgP_p(O��45#���0�;�j��X�?��I3R�|-/	�:��J�Y�T��:ad�H�}d��@� ~�U�"��0�z�N�
p}�XU����x�J��(p��'�6Q���=˩<TXSPvyP�k���x�%�@�d[&��]ͯ�E'�I"�W�{d��՗�����R�'��Q7�����_-��Q]��nüĆ��f�
۝�Ӯz��:'�F=��t�Y�:Vn���h�Pa��	�Q�۾ާ�y�t�%����V��=$���QeQ#��9������薃�(��l�A^�Xl�z�+�;�c�~����Q�odaS�8@�)�8��`%j8�(�"Ga ���/��9��u�O��r�N����z��[hm�p����u��)&S����D�?��&�f��G�3wm��IyPg�^']�p�#9����`��e��-|��/W�(��7Y�_/�����]k�N��(�Rȗ�Q��塹[�~�{� _xv��Ѝ�Ua�:����I{S[�c�aUk�N*�a��"c�^��=���H�y�-?;�d�3�B^�0ʔs�5��C"�|�5LdB�T��'W�k����T��z�Mg)PҌ�L�O?����.tC$}�#�:�������[�&��I�)3��
���l�F��������m�l;w�,�.X�XqH�K�-zM��?�.f����ŏ��.�|�8]�֥��SԪ��:�~�R��a��� ��L�4�3�&�=�EZ��Zv�m�i �0ܯ��)��D�{M���l�wz��o{���@�I�z�t:rI^�	i�	�2�Ц�̙ѽ`a��N2��X��z�$�Vp<�l��哆:R���]�O�-�(^�D�|�#Z7]:b��;P֟�!p���1Y��#���C��"o0�tpr�X���p�}�.ZZ���&I��D�I0�3��gs��Y��"|v���)6���6N�]�Ji�����X��+�LD��ND]�4�4��r5T�G#�W���a�OYLd-������l~��ܗ�{�q�੖=�ո4@-1[��c����v`�W���u`f��z�4���k�LJ��u�] 
_�c;l+GZܹK���	=+F��㣏�Mǀgcj;�R��:7�E�j��/���/�{L;�ҽ�>����`܀���`&Isn!�J�Ɓ�[�$�<uL��Ǆ�8��&g���%��/�fP�z(R�����/�l
���F��J��P�="��`(z��C��^� ��x��8X�+xpD�,����9�e
y��5�� "
�1��M*�����'s���D����c>�����*�f����'�(YO[C�֧RZ��}q�Y������_A*��5�!'a<��m���%\6�)����'Iu����k2_q�l�Kyu4��ew��U"M�zH=# ����m������l?��u�?�|�
��b��Ǔ	��=K@�0�h����~���d0���vF4�]���z�񀹸�w��F��'	-��{e%�s_6nʞ�S�A�q�[�n��k�|S�ҹK��w��鲫n��x#�`T@6�h>\�&���%�~@1N}ᐕVc�K�A�����1%�$Ͳ���]���x�PB�1�b�Cj�!!k���0C�u:����y�j����Yld{��;�qߑ������_lՖ��n䡇V�������(�H�͈,�[�u�]P3�B�1]β�Ng��Ƭ��¦���^G�F.��s�2�L�b�t�ˌw=���;��SPF��u:�<���o�4e��ڤJ���2Eyq��w�M��?�
��������.����f乨K��c��:ŕu�#��2��/�$���X���Ynj�B��ˉ��tY�TH��9}>̻>��Ԃ7���;�\����ҁ�f\��XH��['�7H��[
��Qo*��^`GE��/�����?��wS�-0���U�!�)ׅ��>�2�������B�ه�{��Ï�s棌�o�wx�ܸw�T'^���뱩�O+�4�;TI�}�S�`��]�@	An���vd�76bA����y1�Zԁ#-H���H�Nty�lmdhm�zrq���zk�dP�|��w �z��*5=Y�Q��Kַ��b�b��g� {�7nP��-��E�ƭ�qq�e ����0�P-ޘ9��S�cz�i��7��0�'�t~x�	���kН��Rax�@��4�(�+���9�x��zڮEp^����V��m�R.������\&�wq��-X�>�m�z���k�-��\bL)�%��V���@� /�8t�y�:��-����3P�q2λ�{3�v";&���>�;"|R�v'����^��VW=��!��˛��;qn@͜
�����ǹ"X=2��E����$j��B����|�]�"j�m�M��0(r�<�Ą��^>�q��z"���� ���Y���FT��$���f���p��%�tS��L�YR������u�*�oa���-7^�^�v�4�j�	n&\:��Ck��q��(��=��*�%����>5'����X&#�v7��ڐmV�������ȍޠp�p�(���,�~�ǐ ��F&��T��|n_��������o@��-tT��9�H�v�E�-,OX���.�:tw�;k�$,hI�Xx�^�/:��K�)��݅�f�>�2�!�N1*fL��.���xsi�����47Tv���� �������o��75l��nw(.�O�f���J���P�@�]בk(H���9ǘ\���W,{��I8���k��,ƙ&��$ʷ�������[x_�J%`x8`I���ْ~ƚ%䷞l�a��4���r���Ơk�	m�R��:����'@:���ТQĮL"S��glHI����;����ה��������^dk���qg@E�+�"�[�q�F?��߯�"MP��K�9�S�,KoS6�l���
���J��_/�Ծ%�fI�0��(���1�-����l������ �!��CO�~�+���J�����2�7�{�/y�">R6�����?S4�pas\�d�=b3!P3�]�lZ�Y1k����Z��J_���3ŖbGĔhz@{�����
a��Fpۂ������+t�3��pUC$��.��Y�g�s##�x H�~5����Q R��&ǎE���:�ؠ|�t��!�>�b9|��TFb��{�ܯ�js�#�;!$�)b�q�9�����z)!���O��"���=@d��/.
��&'ϰL˔�MK|�>I��K>O|v�,x}��9Dw`)����!ڎ׉�_<{L��@�d�k��P׏J{�ާ��F<�ߧ��h�MV���U��D��9� �<���������jY�H�������uP��!w�ďz���~�f���̲�-�\�g�������j(1Pg����QLhk��5���Y�ֵM�5���Ő��_h�ַ.���U˖�V��(fg�}�����!���������t���t���|s�ި��U�����gy`��/S��\}�*܈��g��J�U�z[U�F�x	�Һ�ԫD��S�Q��NOX}[����O�I�1�Š4�Īx�pȻ��B�;�ZC�����,c&�hu�����œ>�V�5'�sCJ.�j��R�ՠ��f����w'
�Z@]sUeZ_������mʵ���~>���H�~%�b��D���5�ʇ��as��%f/S����M����5�CS�m�x�P�@�ʎ�$�U?���A�~8����f����G�c	�b�m��Ǵ����1�g�N͘`F��;5�Vf�Ց�[Bۃ+�<�����Ј�z�3G4Ibɡ�d� b�*�����\��t_���ȶѫl���.�,Z�>O�����]Cb��m>��ևt��l؈c *��{��Ł5f���ҵ��e�Z���-�%'�8)��R�O��W�B����,8�dMy��Z������Io��/���úe����O�mi:�x�][n�f!�~Ix�y؊9�][��<��^kZ>~L\�>�I��v�ġ{�Dp�՚n�;uQ���_�-(�Y�1�����v�{]���u�}���n�����?�qB/�|����I��3�ؽ̉@o�T"�o&�L)ר|�(_�ho"j�] :����;��Q�u0��5���xJ{�v�Y�AΗV��$��1՟��Qq�\7�aZ$�}�g��!�U���'���V��:�s���z�$�}�?W����殒m��h�p�Xnע�������9�&<n��lR_�_��0���7�0[ƙi��G��X��� �@�VN��=Ґ�W��8P�Ӭ��~C�&B)^V}����u�a^KD�����
~U0�1q_���b7� �'9�PD8��v]��<E�,M�YR+(�E�o��6n���k�Ţ;�3Gn7��5�oJ@2F�~�(��𯬃8��k���"�������;��J."~�G�Lj�OXjJo�g$�o������p��W2r���9��������l�#�%dڜ���\h��(0"+A��]F�M����J5�zQ�b��[��j�n���	6S�gPzv>��i��Ga�w��m,j��h���SC��a��vLҋ���"���p1N��^jB���|��R6�@&̫o���
�R�Ck�1A�
�h�n�J�4||ͦe>��M�]F;Q*��w<C��	M7��1�����ԙ2��S���bH�R	��$Z�|�p����7ߊ�V�݈�� �uIKlK&Q���<�9~R�x3vm�g�?����5�,�}f���!$�h��^�?�А�'ۋ�lK��G�Ç��W���_��N�RU=��E�V�Tz�TW��ӌ�>�
2�੢Çt3P�L0���	��Hǧq�@��|k�U��}��e� %�dx�7�E�����}��b�����C��O�Y�
�E+W砧[�~Eш�6�`=�����Ua��8ju� ����� G��6��;��DB��w��W����w3��p�!F�^�r#)��.��2\�˱K��d`ttK��t��3RatzO�_ItqB�L�EU���� �Ή�+��)�5��(:]n���q�nh7��Y(�уM��K�@L;���%,��*�E��VN�Rֹ�[^��	^ѹq�3�C,��l`��|8��K�V�;�x������+�h@���������W��_�J5�n�&���!����A��V� �-<�}Fޖ|+�m�0�g�яl) ����R�^�8`�a���Y�.�ܻԜ~g�k��D ��H��}����"�R��B�&D�q5IV��W�L�2 �G����N(,B�jx��L�Y�Q�e���R5���d�r3(�X@
s�&�T+��,H�!�H9G�|(�Dwl�����h���,���B0���a�t ~��-gຐIM~i��Jq��?]�%�0�����Z�vgݒN�2�DA?��a3>�gOf�F��~� � �3L��#��[�LSU-I��,�#���TT�^����TD���"�M<+�%u��~	��fԯ�ݾQ�1�*��]���ȝs�8��0��W�~yl�+$��4cV��Y���ǫ�������S�ǡWH\����kEz?�7����_�����Uqzʴ�������* Y�E��[�/�^0�?�Y�1�����^FrLR!�)�'��r8;
逻s�ٜ�%��b�3O�$wO����Sj��p։�ߡDZ�'20>/c��ء�Ld�}5yZ�g������x	~�1/�VJ�'x/����]l3ɑ���c�>B�y\���cH?������ῢ���V�+�x�;�&O�T�7��ѡ�N�B�r������V0)A3D�v�Z��Q�g��T(��6j��u��	�QL�m���"C>���i�r�_�����n�O*���V�vы�>�hp���ۓ�����6��V4�����zc�C ]ˑlq�j� ����D��{��l�py#v)�������������3��N�X=p-1�H�	�BNB����z��c�@�U������C�����֢�:.%)�.kA�ā���<�5��!�,h?J>2)퍯���<�����|����?���)^� ����P 1�"ϊC���c^\v.EZ�u�"T�ql�fBk���j��B&���%�B��R*f��/�!���g�g)���1�������t.�W$��3�=9���~����l�7�����P)��edj8qf2^y�X��Zςrf�)B&Xr�Cmڀ�{��*�W���w3Ac����9q�B�X���W�l�g�^��m���B�DvK�Hh�u,=�D�_�������Mø�b�E3^e%x$���M�.��X��!;qM�"wZ��=o�F�da�Lc�xU�Zr��Nv����z��v�)$(���c�,_toB!n�kB`)CDR%6ə���'Kh���3�c�W���Vl��}�NX�h��.#�����H�����Njd�I���L�O�-�i&اȱ�!���#� �x���DƮ�)a4	w}�c���*��ھvd��PquH��c���lxKDw\��8DHB(�E��j;9.C�dJ��h$�8���5L��鍬^r��ʡ�7Oe��)�F����:��� ����0+���mgLI�"����NB�A�`�,�ci�SGrk/���lEJN�t���%8�H���U���Tߔ�����4&�=�{�k]��>|NtI�6�1�G���8�eI���a��T 	�3c��%�����,��ގ��1�n�́��.�M�*��f~N~ĵ@T���C9���ik��N��ѴX$q[lD#*�u�hB4?ܸ��HҀ�Xv���������	��f�l���T��M�է���7�7�;C�/��R�����o���į��Zh�1��$e��۹���'>��iª��y�H��  Bo� N�-kEU�8�:㳧����\�Gh�n����؎��3I�����4�xV�,�D�*�dLYDO\��!���};��7����|œ�l
a�W�q����z��2�K��'�$b�r�㴀����l2D+ɔ�'��k�����$(h���sH=il�'��J-�c��Iȅ��ZR9��(׭�f��{��V\c#z<�Ȧ��	�/�o�fCtm�+�@������ �ٮEt=�T@���;�V��	�7�� (��	���iR>�#�Ir�:|8C��?ۿr�}G�8܌u�k1�����З�-�9�le7���H� ����祛�}�v���P!+�L�@EЂqf�~vҀ���H~�| �y*cݤ#���
^�=���i�<zd.��x��ϗK��{��ѕ�g�it6�<�!�<�����x�n�hݺ�n�����s�*���c���T ]�欑 q��~�i<L��g2(�����]��%X����/WIb,�ا�f꧔���e��a�:��x.3]�q 2g��>���)�E�J��W��g!u]�����:�='n\i�H�A.1g��4�S��c����F���.FSB؆��s�2���	�����!���ک��~A0�@����W'��Ώ_1��������T�N��#Ï2$��0�ٿw��Ĥ0s�ƴ�!����`	����˱NO�h�Sj���p�>J�i	8䷨�?5F�J�4�I�=�(kФ3�\iq�Э�KC�xX�ĝ�qFg���F���A��i[�~]Xb>�%ʢ�=�&��υ��Jჷq�~�D���oVʽJ��2��E���M��LxA"�J��%��s�=��B%�5;Da�sM�M/營�u���S��B.͛��k�s�][���k������٤��O��D6H�k�<��6���Aez1��K��g]�����ھ|�����ED��������n���}�Uw�}��{�ҊO�B�H����+f7�x�������[��>.���|��Q(`�-�Xpt`ȁ�}[��pǪ�^՝N$�|�8lҠ�<E�E�F�܀�,��]��"h�&��l7W6q0�zܦ��0���*��`�k�5d	�N�>��A�V�6q�G��LTZ7��u\�u'+��[�z;>��3�CV�,%/��g�4��~�o���C{Ϥ��Y� LL*��P���A�/�����R�P��#}0c�n��!s��_İ�c�r ����m}x0��G�om: ��n����)�ڜ9xM�{�N8�(�5nݎ4�
���e��~�DQ,���倿ԡ�C)V�J9�=gp}�!&�#�q���v4�#�UƯ/�ע ��j>qbRh��J��e)����3�`�}�A���S!R�q-�����ټr����z|~��EN��q�K��J W���B�:C�O�<���1��R\a�V��,jb�L[�#��HV���+"���Nb(��'U]���6Ɍ��&��W̸�j��!�����
h0�#��eѹd��8��*l���O�og�!��0��d��B�)
��(mO��������.�4�|��JJ��c�A���2���-M�@-|���;������Pa-D�� ���KQ9�-�D���G�6C���I�e��w�$�)��jZ����j,�4��$MP�lx�a<��ս���N�,
A�!��x �eG^寱��7yDF"����y�*�W�'Mj8��] �J����?�6B
��]]�w��
��D�]t6�˹gco��+�'-��tu�
�ږ�뵧4�ǥ����Ð�X�����|AZ}��w6�R�ɕ��a�Ǜh
U�)��p���-*���1�5�xk��G�@�6�/�Ὓ��QĈ7I��׎n%��ڄ2(XsbŦ�:%��A�;��"+tԻg!I,�Z3wi��,�y��ݭ��l��ʻ�HGpR�ߜ��$U�гw5�A?�äێ$J	5���j�Cd�~�yn❏am��
�c	;�͎}.��N����&z[i�*$� �>�AJ� �6O+_�?���U53PD���0=�Cqg��}񯙵E%15��4	{�c;�Eϻ	��)��U{MKs��j$��ܲ"T��GZ�
W�Ir ����h�j��T��*m�F�������D��Ts0^(t��k�y�tA���&���w��]7;[+���C�䡡�ӂ<7���]Ҥn��&܎��`5<�l��#Gq��&���b�z� 0����po[�n�Q�⟅C�:�T�[��>�
��\�_��=r��|�)bm��RZ��M��c�A������8�Av�*�:�)��Z��D�`��k��'�`�2�a&ү���d@G@_�ˈt"�z�e�3(���51���I=γ*�l�;c�v�4)��BQ̮=-�7��&�&GS��47�^w�ʲ랧��p+��1p���m���".ho�����b0h�d/�-���i����G!9�=1���z��_�=�����kfD���d�1�7�U�yy��o�qL	V.�b#h�&
�B���pf�8ul*�;��йM����z�%�*�����(p	�1*��� uAao
�y˘�1s|#hP(��v���{�v��Ic���hVX�����Pwg@�5a��Hʾk�%,3Ѷ:�l���w���>t��#Z������ZM	+2n�GG�&�16���n�T9@`b��XiF�˥P�K�(R�Qf���h���g�}�-���bг�H�9P��>���3��닷�H�2��ՒV���z��<�e�_�����x^^�� �VV���(� �X��~Q���rn�Tx!� ����0��o��
�i���iF��y�mp�Xf��r;(Cw���1U>CٶÄ����E�|
.G
,T����n�;�'�L:"�S"Iq�ʃ��5���Z]s��SE1s�砚F���8�~M=��4^4h#����	��Q�Y���<�V�P&caߧ��]PI�ne?y��l�8����}c�aޔMM�R؝��G�8T�AېiW��ىEN4vQq�G�SV#.���Edf�[M.��4�,`پ�{H_T=����`��/��L����w/�z�ZC���l�6�:	�oT
��T�㖝��_��l�u��|��Z2ǝˋ�7P����(ρT�@I�m�p�����#�X2sr����mS�Q&�/�0jFN�����4�dMT.�o��d�5� ¥����a��5�nW�3L��bEq�����<��s�kYv~N�s���i'�����Wzi�*b�1�]���<F{y݃gJܕ�g����}I��� VHiw'2]&�4�S��0�|Ot"�i}����{	=�YŢ�,��=��'��gW�@)���<� l��Xm�Q�Ƀ��lC&�ּ��ZZ���*��P�5
BBdQ�)i����c�� ,�r3��k-ie���ⷛ�$~0L�&�&��w4�޻W]�����s�?���22����(��!�*�aK[խ������Q�/ɇy��3�> N�raGdfOi�PD��~>=t��kcN� B��9������onv����X��,D5rW���+�\�"�FT4��%�|[X��r����U��"�I:�)�js�Lx}r��IUg��o#E���F�@?�wsDNm<�e�DL��-�+�0��r�d5W��z�� �6�A�*�?��Ԩ��g�������j}Ǿc���T�3]�\Xx�MUK��``(��u^�D�S���E�6��F[ f���Y��9<R!Tk��A�
�B�lBRa��d�#i �#�U��lĀ��F򡓸��K/|�sY��x����l���]����^h0��E��c�����r���^q�z�m�?�?<��$�զ>��_!�������Ni$��{X6��b���w�g&����&�f� ���:����;�K�@�����VWC_	d%0�S4]���*�{jfh^{��A�����n:G����?:Ti�KO7a����Ni���L��l�JI��e����p�r����hNBǼ��=�q)X45࿓�e 4�v�@���G�젋xR��>�y��*�E9�t��醘3Dq���۸l9
����iX�Ϡ)�����c�Is����~���@����@�)�&�d�}W�j��H�)���	�Q2�uOg�<�[|D3<a�t �`�&�l [X�����g��lL�Y�9�C���U�iܬn�R,���BL���6R�(�C��4�z�]�Xˈ���L6�]	=�z�*D����I댖=)�("'�Ԧ�0���~K�"a[ީ�wd��^e����y��R��qk����Gg�����;����e��6ȟH
���o�K;�ӗ`���t{Aטp0�'PIl~a����M���ލ�6n�y�)�?*�[*C�$���su�?�(�.�)7
).wW��"W;�A��(Bj�k��P9�"�b�uu䏌`%��ѧ� #(��nJ�z#��f8�P�IM� �[b�S��nr��n���6�BDq�/��Q����-���C"��o���4�2����/n�X���<ϡ��V�f	6i:ƿ�o������S+�(Z���88輻����ݶ�&-հM��;����ʮ�&r�W��:������U�����wS��q�W�?}�������Gэ�,�H/��=Spߤ<'@��/[M�c�f_�T�<�>F�d�(�	K鋋_G���O�S�R�ؽ�n����L/N�m�z XuL֑j�2�5�ۦ��ǅ�h ُ�;�:�dߔ��.(�/���M�1i.,�l��O�c��J����p��v��I�ƣ4������ܻR�Pe���}���Et!��a���Yy{,�"y L�-�y�R��K��U���:�;�,�Ge�ى!��o�bUpĎ�7�/�)�X~��g�gҽ��4v���З��gC�l
 �J)��3���ak>0
���klo�36��������[����'�&�p�̎���wA7�kk�]\��L�e�ԸmYp��/M�ٕ���t�+�����&v�1����M�!_(�&��[�d�KZoe��1�GJ��k=E��l�}7��CI#z��>���B��<��!�N:���P13$���7�ᦹ�=hڼ��NFS˽��À/O�ݻ!�m#_�b�F����0��X��j�F��c7�J\e�J��eo]7s���:����K��T����%v5�)��h�#��9�r�z�#����
ď�F�m�1�_c�w��3�� �w��
L�m���NPX�
R�WuD ��?���g;q�����ͅ���������_��ee�\3E���!!�I2�O���q5��s��%��E�f�G^���j����[l�."P/�!��м\��y�I\�78Rq?��ӕ/t)�`��جXq���H����ɩ���̪�>�h��F@�;a�y��QTuQ�ױ�u�2S|̾V���x���_,��;�Q���R��#&�}.Qx�
��g`��	��w���� �KM��;R�����(<���Hma�����a��HDd�L�0�`/����@0��~)�YO�_Y���iU%��fj�Y�(�i� C1��9�v���4{頪���������с ��\�aōݷ7��\�e2+Oc�Y9��Ko,E��� ��j@k��Z"�r��z�{��A� }ZZ��I���$�V���I�!��j���Y��Z� �����|c�7�0e/�$9��w��Yّ׳ir��V�%<^�2��T���Sb�t��h��z+�s�����/����iI$*�\)l���d��xR2J��A�u��l��Z/�-ª�n�5@�wL���&Mpf�i���G�����=��6�� c5����\L������/݀#�&�k���d�i�wGjݯ7�2����1~�6۟��z�
OM4c��U��^Rq]i�Ǎc{x��XQ=�w`m��-J�l؉B|TQkϡ�	Wտ� 
��y��fp�M�+�&/~t�C~'� �~��b�യFtkc�2f�a��ھ��J����)�VgBӆ����[��$RD�ʉ���rc��\�7E�Y\��9D_Nn��F�K`�	lԝ����8 ��@��u1�d<���'�e�$��NPIrGx�׽�Ҹ,�����a8���ec���Q@:š�LT�
�8�*Z��N�=~f:�a�m��\Ûn���=~Z�#��RY�~�ͅ'���j��&���'�p�MG��wL��~L�]���@�Cp���t*y!�B%����FEon�ns�	Yf|�u�.����[��y�m% �A����*eN���u��Iܥ�T����lx���YSx�u엷�,��Wj�TP#[�|sy&d����`Ж6
��f}.t���>[z9ܘ�*�K�Y�sv�V��l�V��ޞ%����ʠ��?��kK��=^'��T;��k���k�陣~���3�˰��58_P��z�g��S:Q��<Ob�_�*�j�f+��)�K��Ը�F�q�8SN�_ڹ����ur���,�)S��wi�r���E�<#�>A��%�.}�+Y�H���λ�`�z?�ͬ��3B�}����`�ˉe��Fɿ^֔ch'[t��Q�zڪ��[Ė���)�yE�ҥ�,��b��X2�@�����oD��=h�j��� bd���	��z�s)�s�ľV����PuSdÆ]���^����M��HXH�V��̈��/E���x�o:�;���Q��U8	�`ZG\E�C��M$����	�3;�V1tJ`d(�;;u���uB�1��?���:y����Ь}Y����˞f�ֻ�FSǒ��Z���͖8��;�ڟ��̱��RG$˞r��͠ ��rq�2���R'/�O�c���`QȀ���������D�t0��M����L�{%�/���� �����ÆN�ϝ|F �%t�Z�;���(��v:���)��>� �s�B|�??��be5���6������C|?��i���Aw���#�=��G���0�τ�&�
�|-ex�/��n��쀺P���һ�;�ì�������R ݑ���B�!"T8�]Fz'�X��ճ����k��i�	c���
} ���^���Z�X���,O�[�f�����݆ࡲ[����J(�Ҋ�`&��f�͠=Զ�R����=��t��J!�N)M�cZ��������N�h�.���l�!��� ����E���D�a��Qh��tʰ��n��Zc�J1���	�ʜ�(�������Xb��=i��&}��H_W5!�17�y�U�nN��p��(ن�;�K~��?�o�HA5���6#���T��h_�_P׈�?%m���}l�����ɿ({��id�=�2+K�g�����_gs �N�fsWJ�Чuw�����,fW7�D�Չav�1��Sa�������ߎW��m5��.�k�]f��;Wؿ��{u.���Y�	[�������r�S�=�)GLо_:�U�i`�]�-ۘ�����\��q�ީ�t�V�*���P0���R��0Bϙ��6k�+�4:L}�n�����������Lj�JA���G���D+���GJ-R."�� FtY��TQH���2�Wۋ���HV&����U����^eq��V3ؓ����IAS����;�'Z3��R���M�O�1|��Fڌ&�6e��4�9:^`띴��jH���Y����-��ל�*7N��X��Q��c�p��L,Ms�x
����)�"�����96Q-�ҳy\�N��#��w�������r��{vm=�)���|�1!��2V���
�Y�a(E>�y���}��r?Z��j�B4v���GGY7���u���Ҥ��_�u���2琒�p�n��X��I���+�T�uW�e��X Lܺ���,*��Ok2��߉��N|0l"/b�x���.K�'��j9>�����]ܯ65��i�����,#���&_Wo	��"�3r��ǣe5#T�)$t��9�+�C�N��%2�}���[���T&��9d�=4> �8����-���P��}s6��8	�^���|Y �9�Е�1���{_"�M쩂)ӘO3�hTؓ6ژ��O	��M|⪉e.B�e��)�qH�f��L.�F}!�Ի�M֟��Q�:�P.���q$�C�+;l,�ɐ�������i0��K�[���I��bōC�80�}S
�2�n�i��%`��j��gu��sfNˉ�~�{��Ar����%��}[�_��w2�Vb���02�aH�����'U|.0'�{�����汾^�N7(Iӕ
�@E��V��R��O�� ��A����o�p����g�|gn�-�w6��[H����ft=�JVW6A�Kg�U�G"մ�M>�,Į̙y|�}�c��E��	WdA��4�J��U�ʩWt�P�� �#��C�v�i��>}�{�e� /����byޕ�n����Z�*��h)> z��0�>�C�$J�����`BhWs�!���@���C�ENJ_���Zr�w`��K͈��E�6kOTH0�~����	�]B �af�x�G1�78ԦD�Ő`��X����>�u�wV�a���|���GX`(�d	�AH�+��ޫ���{���1$aeԎ(*;�s[rE"Wy����x���c�D£�ƒf�?��-���9�XK�A����>:�S�4C\���.�Cp�D����;��z-��/�;[s��$	�����e����K��}�?f�ƝY�M4ZO֧$��\#�k���EI�xQ�g��qf���m��By=�ʴT �{`��jN���䰃X� �S�v�]C�ph��+�h��Z���S΂H&f�#��غq�3,�c�E����X;��e��G��.l��2 �g�=fU5v�ڢ�Sp֋���<�Ӑr�%����2��bѱGh�c!���);P����i�b΢gAOGU�*�Pr���J9ҩ9<%�04��}V��J��4�i�Z�H�;:��f~E�r����(��ߋ�mؙ�T��^���!}G9���n�ar/(�nٻ�ʗ���k����d����m)Q��D�^�p����\Ԉ98r�T�)2ܢ=d9b��^`Mm���<��f2]6�
��8�&�i`L��V:�&�0��b=�Ġ\\k�SQb�7:��i�p��6�H���c�o�h��!��^�*b�q�jK�8�*2���D��!Я6���v�ƶ�Z�.�!aC��7�J�D�v�kL�f=壤zqٻ�]���ʆa�Ї���V����U��gFI���@Dx��l$~�g�/���6ɴ��~�s��b���	��cZ3to�~CE�ޛ������,��Y����������;/E���s���3|I�]��V�w������z���ȥV�X$�{�퉈U��L@��f9��:��M	f�s��j�^Q���LaӉ��2�2&�)�Kڷ��+������ʉ/-"SY)w?׋��8Wy@b
�z3kWQt���]��s�l���^�2£oT~����=�:m����z��5����q�0������;;Xгy_�[0+r0�G��w��&�N/z�)�w�r�9�Kob�K@m�N�ut��y��ej��/��o���x��/_rJ*00K�40+w|���R�6E|1��b&n���A# 8=c��߮��u륱�_Ƀ5E�]G����� ��/뎵�����>���hoY��ݷ���1Lb��x�z�R\�(���h��'4� ��`�T��sx�7�+�J:��4T�+��S�y�':5��=Rv=Γ���`��}����R����L"*�ϕ,nRЁ�`r?;Sd�@ݧ��l{		Ju���5Qm"�F��iŤ��;LJ�Y��r?���B;0��3_X�Z��+1�d'գ���l��ݢC�.g�Iy��!���Մ ��	�H����
���M�Q<��hH=\8c��w n���Д�3nR��fq�\�=�H�I�侔g��_�Ѓ���c��hx��9g���a����=�P�V���gDv�S����!�Sm�"Ē��%�->?���u+�8���(j�Ц���'�d@JL�����X�$
��d� �;��$� �ޡ'�x�Q:!,-�Ǿ,#�P��Ւ�&f�U���O��@�gc�7�|c��%��yw�fA c����E~���SUݷ�D�I�m߾��˱�=������Ի�c���x�f��Հ��S0����"׋Lg�{�(��1�Z]��Ԉ�D�bZ��oVŁ��h��=p��BZy�E_���ʯw���O��4�?��Q@�����;z9����5�����м�H�bgj��|������,Ūk���M��o���dj�"/����W�������E^5����/p�4ʱ�UV �p���G$���eV��,w>M�ǕBAD��}ˮ���I����Y^�1�u���b�M�!<�4�s��l��ɉ}ߚ�[<[����ODp��q���<���-�i�hIU@�c�$D�t�_�/WTp�3�܃��'�?��#�w6�S���5FkT�v�]�ZH�B����aZhd�&U�G����㯱#J~,2ݧ��OjO��Dj@4"��f�?�G���6L��-z�_�|1깂�Efصs*6V��'��+,K'��W7��>ܺ�������(Q:�3d��>�?�z��S���չ��cm/�CH��:S�O^
��eatAt���,f�-���zaxv�<�����Z\�n�;:G$Emx'zUpT�2y"�b�����YUd��Y�9~��fN�3#�yT�d��� Z����!�p�@2�'���q�z�+ʭ&v���R�iG�����_D��_�hi'�dՔ*��pz�5]A+�ş�8P6i?|�GD��u��� �Ӎ����n�p����Oh߉���$�����3��#V��^'�cb��K^}��q�0�4�a��!��yw��T�Dl�����Ë�� ���iTȶ���	�/����y>x�6�ʾ�B�<��G^J�;��xdC�|c��)�%�Z��-a������1L?)��G��$�h�]ό&W��]3����}�^{P��MZ��T�7���Ѷ���`�0L3����v|�������h��\-��ȧ���a=��dŷN�iD���L
�:����y�����Zz���}�}�E�~�U��ׂ/퐑Y��/�n�M�_�zT�8��U9�=2��zE+J�7��B%�3�#�c���	;4͝y��}�o�"�M�V���eAL����@�����湫"�
�hԻ�0w-�;	_hgfW�_��r��i���T)˭5�Y�������z�a��%(��?<o�xp�+�Z"�/������[�Y�|�.��d�,}�wI#_�5o�O������穼g��\�;������g(H^%Sw�f��� ���;���ن���i�a�;0�lx/�hiNm��S� wc�������yt�����Ȣ��d.��K�)�1���,2�d�*Ǡ�� �0jf�댠�ń��%&��V�le����ǻ�S�s����Uv�'���m%���_;�&C�RR���Pʜ�_��u�>�BL�A7�����u�O�C'e�_��ɼ����S��,���5W��[�������3���ӽ� �'�M �Y�XZ��V|�ys��w#�]�	���I��L��A~����8)6�������"�uۂ�=H\&J�<���T��98o�W�������}�4Z������JO����?m!��I�N{h)���:<h��em6�Ԓ�B����Bۛ����|�+H� �Ꙁ���k�<���hߧ~���ʺ����ʀ%
]�$��{��ba��3��o�O\x<��#�Ⱥ�4�kׂ*̽�~_���r0wWo�h4���t��A3�z�b��(����3��K�}3���aV�'J�{���g�j�饔����n4�ԫ�!�S-�i��E��� S���l��S"�hdG4�����jD"�ڸh�}��
'�m�L�}����Q��f��P�2q�.Bk�@�<�B|ޚS�=�~��UV�Ϫ��6�e>#�?|�0
*������Eυ��g��0�V��?"�^�2�*G��i�lB����vK��cF'�<E
�t2�,�g�a����dj�%E��4�㶎�\���-�U�ѹ>Ғ��O�k�cJjM����2�C���Qh����=��i�B6����1/ޝ���g�Q�/]�h��_��%��}���sCj<�by��w��]�����'o�{�0P�Ȝ�S����e���N��;2�z�5y\�>]uC"��F��`���j�M�P�n�&��у��#�]��:�+���&�ޔ[R*_���QzQ�᡽q�y��w���r\��a굡"�E�	<��uM�F�.3/bw��P+|�pQ`i��k���JG���M��3,�'�-�c�{��
��	E@���'���������^�^)���l ��ҰeZk;�3,I�խ��oN�]LYZ�E,���?PtC�t"�	Y��8���P�I�����j��3׽�񢲡��Wt��� ~�-4R6Y�3tm�rѓ�ៜ�tw-��������Ƿu����d��fZ�7�Ь<�
��J�5,wD͔�f6>�@����x�:�8�����#�fPAW9�y�\w��ʔ�x Fڼ%�j5����7���t�*���p!�a�F�}.�6�����ȗi.�%o���g�3�^w��0��ѻ'���ry�����[�ٌ�ꎸ���Y�$�M��H~�1�}��w�Ӳ}��z�O��o���Ϟ���۫���aE'��e��
J~W�р����Iv+vCj$c�6?x�'���q�2��1�0����K�����(L�=5a��rA���m�c�F$㴧c��������P� �HV�֤8֘v��b6���t/��n)�f�{�K�.�!������~p�|���]�R���$�bN�K�fD;q��TK�����n�T�g}1Ta?��!)��s���SA�)�K��PCCx0S7ff�s���!m{9��=O�'>D�C�*x�Շ�Y������%e��*+�xT.>MU��d>S�5Y�I���Z<��2]CZ��|��{/A�s��.M�V�-� �"��]
�J�&��H�GH�2*
J]�P�O(��.2l�S�Q���ɯ��=�I��W�B�e!R̴�Y�h�ȧ[�w�f�OO�̅�:�v��n(
c$|+�<G�O�����K�yi�ZY��1V�c�YK�w�SulɘN]���Nيᇤ�KjSH1�w���?i�A�[i��.�XL{b���a���{~���k�^GM�H=���Gn�~*��.94���m7�HW����Qp��� ھY�z����ʵ��>����� �ə�-)�F��b�;S��g(�$�ZiGݑǈ� ���<O�#�����[轉�yYF?_��ڕⒾP'7�"��{������P�<�釜�Y2ڠ26����5hdy��$@�);�M=�A�� ���L�.��#rT;���]����@���ǿ,��犩���vQ8����4q����f�8�!+�	B�B1�(K{C�*΅�A��@�O��?G��av�E@��n�y$�؁�8,N;��,ɑ���e�|� �!9Ux5M@N�c�X��~-��0}Ei�0ګ��r��-M�3')�T�EUg0��%>�P�t�,2�l=GM��W!ቫ|�ԡ5���O�idVqXJ�6��[�7�]e3v�>[B�D7\m�'F�u�gZ��/ĝ��2y�{F;,�d$�j,\ɯH�g���J����8ˋ��x}d:�|��Z��v�O�D@�����d+%$��cl"��Gx�J��NU#n@9<3q��3d�`��N�-�S� ��x�Q�*�q8;�g���=�o�'��Т_L�7.� B�֝�GV�!����ϔ4�� ��ۙ��3��c,��槮E�+]F1�D�ѡ!i����SZ��p������l;���p'�;�#��r�?��zo�/�^/�Zѳ@k陼=���,n�t�ś<&G�8��GK"��q{���s�k�6 �FC\d{;,HE
1�Zh�����3r-�Ɓ��J��w�sϴ: |��:3΢@c�'v�icu�*�m/��+� ��lT�#;�v=�\�%�.�p��� 3� 5�q ����<���o�R�N9�֝ޗu� �C#�zA3��7�@s.ΒTw��@���*�i[
����|�p�~'��ɐ��o�kf�ܙ��~���G4�k��b�xs�I3�m �aO�)��ʬ5,y����&m��~�&J;	r��J�VȈ8�ȤS�H�_���^�5��4/0$��a�:�gV�+&ؚ݄$�iI��XMT�h }�^�"��j��! h��V@ �c5�a8��+\!�9��J,�B�v1�����``��'�΂�x���W>2��Pr�Qu4ES4�/|E�_Qh�#�ܓ���+[�,�su�W���9�D�j��6��hKY�Z'C	��@sj���fDX����V<�s��@9����o@��*:J�3��VS��[��b���a��cޛC�JQZ�e ��8��QS�jF.�~������J��FS�,�t����'	M�=��T����oVG��1h-��8C����I�b�x׷<��IKisxKH[�;�IЛ� nA��h���V���}�a�&��)b�Rd��u�.��{d��J��2=���F�Л��L��]G������l�eȟv��>?��D���^���'Q\�p�
IO� (��5(H(+���\���-��]�5'���Z	��8o�:u�,;{.TJH����ϗd}W*���=N���P x�6U��M�O��8s&T�fX:�Y_a��|��w��O!bg��=���S*����+�c.N�o�&D�I�?Iqz�%��3D�Z�2��b�W:�J���j
���V\�>�?ӯ�3ޗ�,�*��&����/5%g��g�3g�#� �z�1��(}T!1�� �=Ʒ��L0Q8�%���z�ɷ�=�t/s4*v�v�c���oYb~��*�z��*!
k�b$&}�T��6���Fz�	�"�mY:�����;+*��^�����)^���V�p���bM*��7���Ьf�M6��S-��薅e0��?��}A0V�^|`�S-L�vԧ P�ι1��i���H��@��m)����-�wQ�ں����Hj��?[�xvPf�&��#^����V�ƟNu�T	.y5��h�==�A�T������'>ioBўR
�R�*�Qf��/�8>^��'8	��
���`F��_rՃׇL���hY��M%7ȮU��"�p?S�`�ȭ�pW�S���!EΌ��3?�!�W��y�<�\��TB[v;`5��a��"
�TY0AZ�j���w��|����m��[U�c�ڵ�Ç��f�=��HN�Ri<0嘍����$��4P�zn\nl�~KS�T���{+���K�H}�x�O/�0�<�:�l��-m�΅;��z8�F��6�BVu���M�.]̊��hq�-��l�)ϕ�(��'<��N�)_�ƿ�$^9�Th� 8���t���1�m������B_� '��Q>��u�pre��6��0՜!��%႘vM���F�8�G��F�z����"���(����4�=�c�U{N���\
�)�����S���	���r�8��I,%V�y<G�����LA��,�Ǣ������?�Ŝ��� o�<�<�^��2�R�ض�D�I�`m�>WT�Q�z��5r�8�i_��w�/�ې���5�򲙺5��좱]���Z����FCY���z����M*�ep���P"��pKy�I/�]��鎈�18��z�m΂ȾSmD� �h�=����^�̆���DA���r\�ש�)�5͉�lܡ�zA=�����}���'��Q��)�"�R�@e>1�=Y���s{�.k����1�I�}��]R�%/dD(��yqY�'�̙.Mՙ�U�Ɵ��o[�91dEo��p<)���%�~���D�
�'�"���B���V��N���/���|AM$��fP�ĵy��!��Z02ӎ���@�Vt����L2��C�����vQ���\	)
s/f���Ւ_����	�x�}ko�mW��8�&?f����@)V�(���NȚ�k�Ex�Pn�ʼQ**�g+GO#r���#2� (�{=#8q�a����@���/�#��Դ�ǳ��Wcڹ^G9���v�+P� �1Y��V�T֓��5{�*��åB��hc�a�?�򤓍\�Po'i�(�eS��W�l�Z�����jLi+>�W�U~'���� ˕��V�%6���L�F�� ;�����7[�tg��1���ѱ� �/ŐUa�9�F7w�VX,����
HHo{B��Q�0����]��Uua���lA�"w�^fz�k�D`^f���._�~,U��ZJ�����ս8�m��hu�l�v$:�>2 ��Y�Ց���>Q�� ���F���m�in����P�F������T�����vɤ����`:(G�mG�P(���풙�����q����0ť���qzO��UW�,.POI:8ə}���xBXg3h,4}6�X�eCvE<ԁx���
���D"�$8��S��^�S��8=i�#X��uLTV��' B�6�1��9�u��n34�<�г���se�ÆM�zp��\���+�p��v8A����2��}�7F4�p�+vCҢ��&���qr�!!�[노n�ue�֋7uݞ(�U���	�gy�3��w�iE��r��-��e������(.�G�81C�9���
��J!b%	��K�(�l.csE���	jo���?��(��U/b�ʪ�`�k��(��2���[1�#8�L���F
��Ō��������	P<��셗?����@2R�]��$�6��{2�b�� 3�>�0��d?�;��#C|���6ޛt5]�G���0�	q�ReX��/G[��[;�l����3a����?��Y��gU1���PB3t����,�hXȈK @(=S�*}x
^�0?����o!�EQ�Қ�4,3�[g��9,�`|�g.X�ݸn�k�@>m��h��h\�Y����k]W��@DɎ���6!!bD�g�T�v� ���ɤm)�7����M��Х�%M�<f�Do��<��ܺY|��	\�֦��t!�S�ȷA�J��ђ��� ����q�K��2�w�����C���P]��^����ZS?S�"%�r�#�ƕ����0�^��y�mY.he�IC��X��ٞ�ܷnL�}O.�`U
E����G�ǝ��S����}�����A2��?]Oc�?P��$��_����]7m���Wk��k�������4�9Ȑ_�z��{�b�g��)]��S7��̆0C"�4-��f�7ӈP�MEŕ
�>Z�H�Z8L�S}����8��3L	�:;���c?��=U�07�ᅀ��B_=K`��s��0�C�H�ڻ���=�\ԍ0Bֈ�>4xm���b�7EM���sڛL��a���#��S�8���n�c%f.��C��#ŝ��ewژ�H���x}��;�v�A$�tT���[��n^��Kvfw�}�W��.�)�a�DP�2�&q@�ڴR/�1��E�Bd?�����o����Іp����Bh<y�^�1��5Q��pmֳ�%�R�Ф��	���D%��|r���i]�~���"�u��h�������6�}���,�2�J����=���Qڍ�W���Q��8��kY�fI[芭^��x?q��Q�xK~�W���E�G�H�-�f*������H��f؉�|r���O m�>�1}ֽl�����]���Py�7~���w�cM�Xk�4R,�S��U��T� ��5л���V�%���2�ױ6�k'wǻ�e��6k�,/Ot=�`G"�yÏ��Fj�#`�oDg����oi��d��+�M��It�ͫ^�n'���_���������܃��>�wϺ1_�{ڡ?f�����0��?&���ԝؔ����nzC��3s[N�������6_�1�*2d�q����rf�ڧ(��c�\s����^��VK�ȣI���u��E��
�u,uкnؙuf)ՏU�I;��M'�B���f�m�B�(KXQ��f�܉3 !F����.%��dʤ[�*��*�g^�"4�&tٔ���O���ǌ<ʮ�x%{_�U^y��{ד(�Jg����V�q,p��z�,J���m����}�Jvq���EvH\!VTM�U�T�k���1QsC��4�Ε'?�r%��/��4���$�QJ���K��m�B�-լF'<Ɂ�ˑ0�vs��Uy��s ��q��2�8v�3-&��"%�B�s���Y�����K�$�`}�X+���е��փ�=��y��^Y�3H�:���h�+\�4Q��)�w��X�����.Y�"����)��Q���BAO5�E�v���HL�״���Y6ŵH|7`�j[&q�:i�n�,1�e��(L+���9�Zs��.��ˌ��X~4����x�nԟK9p�rѰ��O���.E���{V�'䦟�����R��LC+7?�D�G@���>���wv��2咢~��-3�V���� �q�"�4�x;76kn{���Ҵp>p�b1Vޝ �����s�؉�iyƷ�Vd�k3/��8���^}��o�����̛�uy��3�'�s~J�ʦ��j���Dx��(���G�X��0,9�#�n��'-��?�B��#��5?-�	���s;�r��8#&�=�Ɲ��k��ŌV�jY,����פ��̡c�\~�߆�ibp�i�'�y��,k�����(�S�i���L�����Z/�*Oʺ��}�Uj&�x�A�r��ױuZ����75�?:-9$�E���(!��g~�O�oH����+e�D(�l;�p/����781��Wv��������);�Z+*�M1r�G�\�fKP��(]�LF�c꘭��䑼?����cN��]d����C/{���)���["��/^H����~V�\�ߊ5V�|L�.�[���>�����0ڱ;[i�Iii[��A�z'�m.��lC17��������P�= �Vެi(�p�����{<���\��y�%)�V���h���%ݬ,j����uBp_ὥBB3A����u8ݲ��}�UU���ƪF�ŢV��0]��.���ӛm�S(��X�ϟx)#��J>������H���_����6���]IG�_n���Ds�����x�V0�;{_�C��tc�h���s���[���'̭�$�Gŷ�x:�~~��*jXjz���y����,�Б��5���Q�e��[��
f��v�ʨzč'c\�-5�Վ��-��E����e�G��>�p�6ߡ���%�1Q��x�@�*򶯢]�C��( xc���G�{�ud/������<���|��7K�Nm\�M~��/�Xd�����=X^�X���0��x�@ޯq���k�gPQ��f�N���V���)Oc3�p�ԥ�f�Ʒ~���l�:�l`���������Љ0�mLW.������.R��Ǫ���@̈́)��:�`�?��:���D�AŞ�%1�{U{<%�kE���D�� j���f�\;��\���Z�N��	�`��A~��?X=�Q#��ك���W��F�|�0���$Lu�T���v�C�z�����Q�<���pD3��"�	���ne���w#�OI+�F��4��t�X����(����ʲ,�V'l\s�t**�eĜN�f�'��+?,3�9�[�Vs�$�p�����J����T�[ w��	�Ұ^U�_�5U�"W�Kf��Ԇ�CSY�1�)�&�.�(�O��%�-}J�_
����T�\ل�˨������ь�m?5W����~��{)Bj˞a>���yO���*��y�����7.H���y�
��\3tY�*���v߲ϙP`��M�p�Ec�𖵆1K���S�i���bG�V��o���s�(v󝽣�zOe/��afU� >V����/~�s��!�ؗz���� �q�o���� �� �>��� �}��Y7f޳������G������O�&1s-OF���@j2:(��- �ĳ��EO;����H�JaA����n�2� ���7FjJ����W&�]��]e�H�j���i�Ѱ^�#s���2��<�R]Oo�
��|Y[+��UҒ�8�E��>�p	��&����_��
����R8�i���T���R�\��U%�� �M��ב���oɔ%x�
˶���6}��&BVK�Bw���D�h>,��͟3�9��U��ܥb9U�.�-JwB���z�2R���쨵׺C���qc����E�+��kfeF�����3q�� �	����o�4 e����:�!e����u�����.qޓ{^ ˚P�u~~�v<J��s� �@i�؅�0�Ha����k�oW��O���,���"�݌���fq.,�����(�R��e�ϛDe!M�������;�c�7d��c!�*\;��'{؁�i�o�ō �Y11kW����^ڇ�}�vPP1KY���<N���a��'\�?���Z�ƣ�:i�����09�:;'�|&&�9��|�US �dXv��\V��]�u��w�'���o��3�����6���.(��m�/����c ��ַ >WW�=�!v���Y������~<#SnA�	�p���@n�7�H�c�TKHHn+���m0E�W^`/��sXU��!�O}�U$�x�D�	T&�-y�c��"�*�빬�����$�[8��*x~7����B�d����F3�r��ʝ�Y�Dt��hw���$i���:����A�Fsv �l�M(��L���A�q)�g-&�z62`y1�	&�d<|c��e?q���R	q���'��I�3<�!؀k�2j��N�p�X��os��*����ϗ}i�Ls��i��t�����8õ�$�J ΁�
��!��`�����%��am0®�M}���oT��o�L8��m�q%��h�(�,�c��x�:��&Ua�pHZ]|����1|�ZH�:O��2)�G�G�_�(��l�w�l�k�خ��9�0ْ8U��e��Z�
��]8=�N�[T+*��r�ZM�2��z�\�R�y��J��& �<�2e���*"�M)]J&��N���.~2u���n�=A��D�®�(!U:]>\I���|t�	��D�,����+�NL����e�����K�tv�.��^ܘ����䮶��) ϊ�zmoB�뾎�;zR�"Äb'D���W�.wl���M��+B�Bֶ*� K�n>7�Z���tӰ�tm�P<�*������y1��uT,|��[��S�~Y;��v���`S"�[&��'V9�f�ΙĐ�=��q�ER|AQ�n{�3�d��T<��TF�W�口�)�����4�7�o�bG�F���~8I�X����L����(|'?����KZ�pe�[T��B~�Ќn�tM˛h ~�t#M�Z��u�V��h3�V��s-y�9���/��x��4;��C5'��C.K*���>*������T�	_}d�<L���-��d�s�����9�{Y�+�P��EI�'�瘃�O~��cxq]�Բ%�"�v��#���J=\W��Яn"�f. �8����w��ce쩭�+�s���a,�"�O�Iu���ì��
�*G+���%�իQ�"���y����]'��� �V��"�Bi��������LH���}��Q�Z�I
��OS�N�w;׸�gd�GG��8��tPh�u[_WKbw?�[���Hl��a/�n�q�o1w+r��_��n�ԍ�e�izQ�)3����n�ee����J	�� �i�8ɜ��~�2�^�-�v�#?�w��Ir�\}F�ZQ)�t*'e �3f
�j��~�R�Qs��V��t.ڒ�I칳���1sX9PR��4��u���J˰�TE厧����7VU�z��P%R7��QM����=��$j�a��;��M��g�&��_�����]GfV����h�?��2<��֞Ȕ��{�����{��h:6����;m%�Y���4	��e~FKX�H�u]�
�d���O��EJ��FC/�x9��0:6���5�`�36[?�4��LT���a���M�~u�;��>��w�������H��d� �!�j9�"�B�ThD�Wo��9�$����
t��߲�iS�r�����y�˭�l_�+���@�-a>?I� �f�{FD�c�۶u_7�؈ʆj o��]M�T�-&L��:%wU�@	��/' ��ؤ���M��o�O��XonG��3��8��T�<��d���E�Τ���x���ã���^��p��@.>�Ô��Y�x�Y9�Zy4p�}T<���x��7����=�J� �~f^��@u>@���ſ±�����J'����?�х_h�pV���������8�
��_����V��i[DNVy�����Te��2�{'�M>�ߊ�D��1�x]�$eF����<4?��Vy}��RǊ��s|\���x�\Α���k�k�yx��,޹����Y�bs,�nX���q>�ک��O���	���m��-0x�E"������I2���V�'��)�&��D��GҊR�C����(P�T��~'Z��1/��YG�s������y!�X����2�{��m4E#71wu�ZC���O$+O�|�l)go����.u�~�E��DLf
�� +��m�qރ/3�A�b~{���v��=QH+���Q{�Qp�{ñ�4�i�G�����C��f��ه���
��y�M�Jx���.��J�C�n�|U"�{:�/��z��b+����Γ���|]��6������lh�(x#��Yucg"˥4��k���l���	0P�H��+Bp�({�ps��|]7��}ث����JUg�д�j��"��}ױ��[��T�֟�G�郇����]������rh_��Q]�Ys�2���*-!in��~�:_�(DeZ<U���6�؅@�1�Pu����1����I�-u1Ο�w�1�P��ڽ�}���"���^����k��9s�KX#�V�e�ITw��0c[A�|��͙���?QA0@��P�W��ؤoC����T�z�޷�z��l^Q�7�|Nx��c�/:��@�'� �i�Βb��=�fB"�N�1���h�/�ߦ�I����ƁJ�:�B 	�4%��e�	JKԽ�R�+(�0[9jY�T���� g'�+�����н�z�,����k�oS�쿄i)��;0��j���=����|ʬ� ��s��}�r��<DUH�BnĽlM�-o��r_D�,�V��Ef@N�,�}~:�������5��3�c������vK:>�]�#���b�g#��>e���ko����SD��Bx{�\��君����:�y�( �e6K7�ЏO�Cc�Wc~��:O�ʳ� ���&6s�Uw�Є�����o��V?���r4=�{���;�mWO��,�+z��}�S���܇Il_��M��g����ɼ�9c{Z��}�q���6@�5�t|�%��\�Qo�m�O-�������g�T{3JC����)81���|=�XM6�F�l���rrl�?� }��>/�Z�s��T��JT[7��Q ������
�$x�nAR�/[�� ,]��޶.�@QL�$��H�p�wM}8O���ُ�צ-�R����ׇW|OQ�O'�p���w'�m��SA�:n,�Ѕ@�g7�xSf_F�ތ��We(Ϫv�z�,��� ,�ϭ\8�;�"ލ�mc^Y�?)yB���0�ա�{>�9h������WH��?�b���"I�m�]�?��{�Ƭ,%�I)�"M����R<��N0�z�U*n~��)r-���;�xB�d6�o���%�B����?20�4���������|�Z�2�ӐĪ�iv�ݡ�������j�y&�e`|;f�VT8(2�l�XR�\pm�L�W6^VD�|{����u~�����n��T��ɮ`�[9p�dqb|F �$��\�-+: ��~�~�bw�7=ϢI��Z�S�ltƚuO��L�U7�f5K��g����%�S?5�s����6�ZO(`T���j����.&7��²���/����
��yV�U&�A�K�l~k%2,��$0���g�-?4�Xڽ�3�ŪfI鶛�)"���ե5��n΂�fsT�]�4FW
�?�{A@Ro��z��v{b衰ɟ�/#?�H�Xc�i@Ǥ�����;��w��͵#��U�Db,�~mG9���R�k��Tt����E�/��BK�Ǣ��i�{����E�$ہr����h��T+���$�u-{����i�(3�����L��߯�#�1���z!�-=ڽG\o��������?��q������$��#%{�E�?��I���o��Ǘw����0N��ؗ��- �V��<Rmȯ��H�N�j���3AP��`��/�h��_��p�}�)Kp6�M���m���7k3� ���!m�w�M��wOc� v�����J�� ��0�&��񥦽RZ�Vs��ņ�Ju6��Oo6RXZS>U��6��h�[���E���hd���P#_�+n<L��n���D���@�6��O��Ⱥu��=,��_��T�Y� ��nG"��d~/V��2�x�0�={]bQ����.5f̍Q^ю5))2�IQ��~zm"�g�|�M�"/��,
��j���U_b���p�XB��1@�;��� �}jF6��\u����-��E3�̽�m$������e��eX��w�L�T���0Ib�={����{y7��Gj�#���Yίkʹ"���N}*8�dg�riƸ4�E�=��j�����ǵ�:� `vh�XT�av��iH����*���]Rn��o�x��j�XzO�*�O>���}<��o�y�!�N``#"�vY:��_�1_+��h}A���Vͫş����^�y�h?wӗ�V�&(
�s�����	RZ�z�y.���d�x/P+a`NhZXӋ�u��fA-��N�l ��!{��a1�T����*��3e� '5��R��㷍$�*r�&��-�%Gt?:M��Z!�Sm0�!�P@��9���D'�7�n����&���)N�������Nc'�#�t_n� l���ߠ��%O^Ng��	��%
�J�+/�;���.���c��_Rpx����/=ԇ�4Wkh���n\�1���h��������+����kM�!qx�����L~V�]���Aߢ�L�8�?ԝ@�$W(�s����G�i-b���)|��w���xKQ
�čOsoɚ���6E��!V�����15������C�,S����U��;P�u����
��O:�5I[�@�`@^]�iBP:�><��1>�����+�X���ax�NBf��t}�F���ya x��H]ZDP�v��LV"$�����Vx���H�N���x��|��0� ���u�1�5U@��H�g������-
� `���H��5�?X�� ���kZQ�G�ZC4�*�F��]p��<�h���Z�����fl(3L������|5^>�<Gq�:��8���0x@LI8�L���a F�X{I����+V����W�;��A 19�����ޓ�unKu@��2'eD�=� ��N�X�s�h��%��՛�P��䑌ëܸ�_�M��x�ç�$<VP/�7Y��e��
HT�Sl�()�QJ!c�Tup��A��<gVE.����������p����/�V]�ݥ�C�'�_O�^�d������[ge-M��~�0Y��p�_��߬�(ݝ�:�?N��w �������Y�)��;l��P�m�Y{ڟ�����E7��&�y{�!�y�Uc��.~��ᬵ�̊���%���9��-(�o��u��_���]k��\=��
��-眏��T�=q�ՙ��� �_]����;nIп�J�4�Н�c�:�o)G�2�&ȸ\p��e�΅Y����g�R�bJMR��W7��G��N�� �׼���k�7}.w�t�-�]g�ο�]�%-��k���=����>��F�SX懡J�ZA7�a��ř۽�`X2g����A�p�5���ÞS?�w�<�.R_iH ")����-k��P��d��8fml�����h2���K?��gA#�vj�B�X�S��B�t`G!��Rt!�!S4>�Sp���P�����C���_�NB�l&υ�7�Gq��T���������(�F�����r�������p2a�
H�^��]��a�Q"f~�!�o��=��X;�^��F�Q��s�4�X�_9G��Ad\2�1�� �/6{>�H�5΂mn��Q3	F�Z�"�T���-��P���[9�1G3=��$x��_�k�5����^l:VF�3����EE�tUG��t�i��󵥪��/S�$�r!Aٚ�P��[�;Z�M��ĈIUG��{I:�*"�ә�M<�כ���N��o�ԏ�'��,�F��"} ���?���PkS���L��e�+J����UD�W�%���Rݑ���I7]i*p����������y�+�����\�
�A�0��gw(�0%�t�d�Tp^C�d�M̺w۫�W��f�tZ��١���8��G'ʓ������A�!�ρ����;�I0����|�$�0GP���+�����F��^�Ф���$�z��ƅ)�.�YmYpO���Qd�C%�>��۔�$�cK��zW�'S	.�t��������Cl�\`i���3����p�h�pZ|���폿+oˀE�C�w6c�@d2��^{)}��:��jz�݄��l�5b�4�xQ�?����$ߺ��#ف���-�{I�v.]J(�ٌ��WnUE��A�!r(�+�gv�T���G������ף���a�ë-�}��#��7.�u�*솲��Q/Dcv1��r�9ڂlEq�znWŇ���W�`f
�Y�!Yh���qkfO�^�x��xI�]U��%�0�'�:����F �%C�x�Ƞ�t,ZU�H�����7��F���N|�ݾ�|f�}����r	�vb6K�Z��*=f�nAj>���_�i����U��?��:g>zC2��]�p�2
my,>пS~��}l6Yb�Q2�)o�Ĭ,���,�>W�I3E�C��V�y6>sG̤���I��m���|��z;Pߛ�G;��}S�e�u�~W��e	?�	`x9��~��cI�c����z���ּ���Ѻ�������Т���h��j�S��5U�p<�<R7b��$^׮��n|����/l>�k%{[K���QÞ`��`Ѿul��Hp���y��v�9S�&U���������H�2��~��ʺW�d�,���h����}tj��ӍG�a��?�\Q FJ-H[<�n��Sdɲ^QY�Yw���va����/��u���=��GN���5��~��pځ)���;���.�P�R�2VkO��r;�-�t1�q�g͆Ϙ���x)�b��a8�k���7~R��/�/�1z�.�_�Ĭ�Q:�^��.��y:�ͤk��:o�v���;MK?���{�ߕaPYҺ.w%�/�R�'@-�������=�9"�8�*O^�2}�9԰BLo��jKMT�?|^q�&F c{��m�O=�3N^�l<���BV-=ܸ��3Y<� I'�T+�����HB���P�ZB[1�����|�e����5ݖv�5\n�H8�!Y�A���G��OŠ�r_v��b�^�͡�b��ww��w������6W���$ޱ
������	P?��%.Y����|>�D�շ��ݱ^`. Pn��<IW�ܴ�ss�>g<�~��U����5��]Q-ί	������3�B�Y>�����-�bFG(�}�:~���\�A�l��ǵ�\vtߗ�Ȥ�$X8�,R�Ȓc�-�P��*+)��;��t}�u� ��0uf���=B��aG��Jk��l�zkW���#��?&�����˺����k��L ���[Z�!� >S',(��ۼݭ�5��-
K�+Q�����̑'��W���2F����B	��6�?��3E�q	�V�4�=��I���%룅��S9I��Y��j�Qu�2-� �H�m��Ǡ�AKg��ڧ�:J?���;�'��:��5����{�>G/eG\��tܷ����������O^@
��r&���*|ۋGa��MKP�;C��ץa�d�ۍ�Zˉ��Pz�������$e#���J�w�Ӹ�KWY�
��
˟ܾ���%������~�*�
�Kmz�&��5�u(T���Z��Ȁ�|�4T�������_����3��8�̡F�$�)@nۅ�nj)N�`7=�M��L��K���l��a���&0����]����R;V���8�n���H�X���t�{4��PB�8�H[!!�����5�f<��{�T��R���Ht�!Q��w���Bۺ��u(Ft)��@� �Y�n��0i�������P?J�8S��t�}����B�[z����]CzaO���=G��"qd�yU-�&�Bxl	P�&��{�������MT��&�*��RX%�i���BA�g:a��ǔ����!��63zKh�>���z�Z���j�BW���?(�8�H_������u�j��F�lйz\�t��|�tk����j"��8CT�b~��V��I��^��w�~q6�t1���z�16���]��u|�QKD�v$rK�l�T@��nm���B�2���ĩ�,Z���fׇ�FF~s�E6қ�����&]�"����C������c�My��MW7qQ����*���T�U��C�%�=jpZ��;GҮx���+�'�q��o!�%3�Ս'{;����yu�R��<5wѺ��֡�)ל�C��l��g�K^�>�|� n�W�(ȌK ��K[F�#Pv�( :#���Z�T�`��w�=Tz�S6��sm:Q\t(��PU�k#����5���R��.���}���D)�?����#Qli�H=n�Ͳ'�] $	�8)�*^�Y�����e�0�ryv�),Y0�'�� 1�r�,>,Ǘ+<~���`���Uݐ+�<��~**�
䠋|]�	��
fXG�kWHO�{�x�b������x�|R6-S�Ґ�z7������o��o���k�MN�,�����k�Ҩ2{;�M���`����]��{������y��<9Wn� �LTa����g�.����R�v�W�Z3�d�ӷ���q�Q��">6{�<W�� ܹ�#�sc�g�����X��!�谫�k��-&�~�h������s���i>f�@v���[�&���ɛ��o���j�ǌ��f���fa��id+u�<�����(K ����i��\~���
�u�?{_aJA_�d�:! }F2�6�e�^8D�T8��.мDD�΄'F�/|�F��H9�D�rD���uI��L.m5�O�^e*Il�Gh���o?�Ww]/��5�0�ދDF}�ϧ�f�|�E-\�t��}��s|m�i�}!u݋�ɓ���l��ޤ��K۹Y�>�U|�̂�`�[8�[)��2�;hKU���E��ϴj���C^����o6��)%	��e��R�@�=�o׈��T������lZ��;�"Ψ�+�9C�s�0�j1��X��x���Rn�v!��q/�ofy�H�b`��"�uM��8�)�`�is���$G{��K�ֲ�3�t��k�"���V�YOZ�Ή�|�c� ��6� �%$�*�_�Ml�RʛS�$��b�����r#{�� N�i�{LX�Ï���#�-kݳUxq�ê6��?6.�Y6�vp�>�A"(��v!���� �Z�}v�}��ճ)����;��9����O[��n$\�6�c��O�'/��C���Y�c8��{��F����T^gTI��'���>��j�i���!��ps)����u�w^����GjWlu/>��ЍD�b���,ϗ*��t��t�Xn_R���MlO0������������a��I��v��A������b���yXC/��n�����B�
5�){/���p}!X�a�=ƾJt� ���(�i�^O����O��L�/�%����E6�Y�����R��a	i��8�r��nR�r�k�ɿ�Z��]�gm��e�3~]N#6����*��p�O�JI�-�T���1�N��Hb[^�3Q�h0��y�.�ݨ�+��B��E�siukE4�v���ƍZ7R
�6Q��g����-0��̔�n��_iE2�ۍ�S����.1��3tb��zd係x��M�x�N<�us�������GX�vh@��q�̉�Gͺ��tyȤw�^-�O��Ȗ�&�(�X�3�|H�)�\砍~�Go��y�3���S~���3A��rP'fp�ʓq�1�͆P������Jo�uO�}�B��I?��*9�b�i��#%&���1w�n}��9����,1��z�7̄���M��|IԮ�+��i%��q���ӻe1D��B��n�Fֿ���Լ�FZ���"�nǿӏ��-�ӽ��'߉`J�A�+��4��e�&)�$�l����T&����a_�e�����D����k�$kB��b�^5����8�O�f�
���ʜ�Q+�Hz�$��F�Zе�d5�����#�������Ʊ4d᳁�).�,�<v���BL�KJ*� �MS��k�2��e�9CZ�\�:3��
JR����ϙ����	�e?xՏ4�v%ig2�"S���,g������uM>���(P��$'��
e���X��Ӽ�����>��_-�&�5( �QD���-k[Hݻ?.�^�d�YLk��Q�'�Z�������xf>�:.^��O�e`3�O�|��QJ�lQ���ڟ�`R���s��0�	�`�`���g��F:I�|򊋦UE�.�[���?�>���0�KLXV���^QR�e~��\F���G�X2���jgg��M��;�+��`(:,���Q͜�43���͡�2�gb+C��v�,`��fG�U1�#�+�TGQJ�ѣ�[ܟ�k���s?@Z�}-6��E{ �F�L+�}w�$��U�ZP@n~�դ�4��;e2�J*}�I%]�4����Rv(����e�������&��a�������,�:;;��/ ��Y��2�SǀF�:�4�$n[tH��� �p�!������� �.(Λ�2��y6|9�8Iz����6�jZ;.���������(������b��s ��	e�7����B�:"NB����J!۶�
�D��3�(������k�\M��R�aM9Y��3�=���gҫ�-�b���G��[d�"�1=�m�/��1}t	ԤT�Y�A��Ӭk@�	�N��?�wb�+��aZ��k�J���E�����+����K�P����â�y��!s�r�!���y�\0Q���� ��vE�|-��Hdٳ};moq ��Ѝ�Ɖ{k��+�������
�H`3H����uc$Ջ�"�e��|nz�u<|LB��bF*�&G�μ�i��a��.g%mN��ٱ�B��&}/b�	q�7��0-%�d,��G�ȸNg�L�nwCV2�(����e�T�X�b��)�����ۅ��r�;ETΌ;�J�7�rE4c�Q��qمSvTz����\e��v��ۙxsl(�E�b�Br鶖٠���s��	���*��=��d�c0�k�\L�����C㈏��ħ�ب��Φ2{�ϘHP�,��F��F���3�sX��t���!>���?��ف
���I�x��]�v����s��W4��_��Պ)�G�!&'�!��o����k|>|e�=,��a�*<�4H&M��<ռcFR�0�{*�9'�<��:F�O���6�������������L��5;��/dB���}#���6�]$t��.zn���m�g�#�����Q	����	�N�z�hI�}��-&�`,�,	n��Xb��S�T|�r=,���0ѻz`-MKy�����J&�c�-eRj"��/��!�x���fT�r�{��f+�U N��"m���4��p��=�fg+��Y����4�s�k��TL�q�K�K�x�$6
�zM�"Í���� �G%x&��=��K�L'V�Я#/��n���5��,(��{�É7�='2ҌYQ�Z�ہZ��V��4�"�+I{g����I& OIL��41��=I���D~�k��Ŷ��?���t��h`\I�	��k�T��q�ֵ���uVEI<%K����t:�i�jΘ���r��9�҇u� ��H%���y%��Io}ݨM;wk�#ԑED&��[`�����)�p`��\Y�w>k���r�T\|�{+DXD\н�&%޴eq�\�..;�$���ꊅ3��\�#�t�M�M��I3h����ܮtP�\F�X0+<y.����P{���_%��ʈ'��l�C9���:�V�G�|�g��-��,M����*Q?��n�	�f�D$��[;��:�w��j|Ap�JO����z�t���:7DJ6���aKƟ��Q�/Ͳ�*��D�Iwj��!-LxD.�)���7;��}�M{&r3T̬Bb��{?�ؐ��eby�t������5�������»F��KU�^�$���-3����njS ���yD�����߇JaP)O�2�arw�p��ݙ��p���m�xa⬙�c�B�~,��e�b,�]ի�6`��w��pՖ����_�\�)Y���"�5���~��9�,"K�)c8Ȫ8� ��<8kd�-�F'6`������M�ƽ�Y.�h4�� �k�0'�o���4(�;�L���JV8XM�xmtjTX�;���,�E�*��39�g�|K�qY����JQ��"�dt�9 �}3�:�z�=�`|�'�q��W�6DS�	U�\��:h���l���m�u/F�JIq�06c	�ᶱ��� ��h	M섿�-e;�Y���8�C�/4�FI�^#�v ۢ߳Zg1�<��/��XE��}rSH0�7�ߚ�F_��Y�*��w�X�����K��|Bp�p3����e�|_�ÿzk̗��@J��G�M�f�iB,�`�ZFsM�q�p�T3sQ��%e�W��
)wb!�*���%�3$����M��dؾ,)�(�5}r8�l���f4��Jo�]����l�eΒ��?����@EJ�M�M@���R1m�'X�ك����d�C�0�Bj?f� �@��1׈y�v��Y�۪H��sE==!���Ve�/�f�5�DI��R����V��qiO9}4���є�p�ۢ���|�m�����P�w}iKp��낌�܀���GS��M�,�{h�I�� ���!R�u%p՟Ϭ�d
�3K;�ŕ�"���Z�Er=dGP�vf��fu�EƖo9Q=�W���ra�A9jUǹ˃�M,x��f�����v��5�T��w�:���kL+���{3ɐqQ�l�z�	ݕ�.�:�8����dn8β�E�/��ί�mbc|���#]My[&��gq�(�w6B=�.���Bd�C!�u��^��r���.��~����Pw%[�kZ�a��l����]�j�B��$�-�.'�5ie�jT��e~�ρQ��J,R+sa�lB�U��9:�O�[G8h�S9��o��lf^� xմӆ8�ۇ"�"���ԮU7S��p�o������\�3�ur�66���l�z�y]�ܸ;9�u���}1`_D�<SMcc�݆б'_�1�Y7�v�`��rf�o���X���˷�.7�@BC��D���y_Ҏ�5�5��2��{�AN�j�QA�N�S�aH��Nf��Fq�a!���K�C͔Q�VD)�?}���͠���C��T�cŲ0�ـ_�%�ؓ�eZOr��u[>�c����fC���f��=�qтZQ1��*�\��T7L�č`�o���GQ�h��l�/�<��j�Ib��Y�־��MHH���%+��~������		��8�O�H@a��aWtuڵӞ��N��Ĩc^�'��˫�����f�߁N�ك]��
�0�R�!�o3�Zme�%�!�%�Ί�u�$�h����.]������.<�[��;!��tIQ��^�`ܟc�4��:i�#l��_��~3�0V5�fB�A���
�<ȿ.�*Չ���1��*��J��˹,�����!<�d����5��	��zxv0ŅR����@��~��Sa\ɖ;�����E���:��[զ��g[33��I^s+��w�+��\:�
>2a������̏�q��[�^������?2!(VN��Er�u��w��0���5:��:����>8��p�T�=v4��Pˆ�T �c�hUh$ӽ*J���5�SP�U��wbO���dS��j�n|s]z��1`�۲���]��	z��XiO�8.럝龺<���5��I�YOq���|��Q�D�b�ˀLj����Ir.�;t��?���)a���T�N'(. �Wq����d���h���.�
�g�8�>���ʼ����O�**���3[~C:-�{d?�B�m<����
J�13%�w;[��[���8��l�yg�2uߝ3@io*���!l�L�����=���Ϸ�L����i�L$DA��b��K*F��n���b/J�Q�`[�U�.|oUE���u���C�Q�	p����LF����xn=�'<�ط!a��!�v�H�@)<_Bf���ə�|2hm%ǕSwלH��|��~OI����*��x��zVZ+	�4|��A/K_B� f�ve��%7��P�*J���9��lb@��Ͻ���Rt���4�pկ�笠�V�\�H�R�Ub�D�.xM�1�[�[m]N��`�2�gl(�c�Dp��sԲ�8I�4�������ސ�P'aU�E^YJ��1�T&bp�:���V��9�S��)z0�b��s�g� `+SiA�9ߦ��)�;��^Q�(������K���ȫ�x��.v)�ꀒ�O�'�Ѝk�YyPC�+�֟*�|�9��g��7Ϸ��?Q!Z0id�=������v�ѹ󾽁�M�;�w��<�
S%^��/$L�8������M�n>�yU�33�Z�������"�SF� ��I��mM�_+Y��L�zǡ�Q��8�`�	�UEz]	e�� l���\����x$�Ɋ1Z�3�<���n�����T4�m�����%����3a�d;G�T�3����w���oQ�>�sW;F՜����F�}�=
t�/�x'��H}_iy?zu�Q�In�*�m��L�� Y4�G��ד��*�G���R�)~U������PbN�BG�^0UGS�ì֛�*26�ߪ�}>$�}�0C��J%��5�ݏ"�Q�Ìw��ʭ�*N�t�ScȔ�F�^C���-�g�:#��
��ئ�����f?`Y��8EG}��>��v�
�ʰ"ͬ����8��6��E��U.A����'�%û]�9N:]յ�̚����뺞V�`�`r;m�@0�'W/6��oB}�&��7�qǏ
"E州�A>R1�2�i����T�Z�i(�%Q��yN�}k�׾
��F��ȥ!d�5u��4��kGHp)���x�p��Mm�R����T��V��=8j����K�����Nr9'�Ӕ<�2�����mH���ە�d�8Ͷb�xtv�;�H�:��n�W뭏H(�]�R�e�y��Sw���`Ҳl�g�ʤ���A��Z�~n0�sӢ�?2�����{u�&4�\;����YE�����'��J��Y��aA�Gq��BM'Q "
*���j�S�w�&9�!�v��'h�g�f������t�JV�7�����w�֚V��h�/goF��E�;$�5�$�Z�Lw*zrZfg�e��+�v+�x .����Z�Ji��T�O~�f���A	���oX ��Ɋ�j'�|����<�=�W��R��r_h�V}��q�tVP��d��T'ð7�v��΢
�i=�al���8�?���-E-;�r�C�G��=նyR�@�c=Ag�y����P�wo0dx���?�����;28��x��u2U���$�*L�8=˚���n����n��a��x&�f�"��ca�}���qiN�W�K���_L|�
cꆗ�-D�
��P�׶�KÛ0��N���l�%
��2���e3_ke�\�m���VF�:�H�K������>�����1+�}�'��f�5��Җ��[�#�h�k�D�q��
a�3Q��=B�s�����Wlp��V�<�}4�H6�Tem���5���ҤoY,��ୡ�_�6Y>���Ț�ש��i�V�S�p��@',�Ԉ.�R_����wߒg���y�^g�3n�~E�/����MpG����kV�Y����b]?R+���ie�5��"Ǭa���F�)���/��MO!��?�UӰU�,��� �B �B|��M��lkO}��<���<ֹ��v�t�44�>xb�	Mvtx_���i*�#/�ҋMu�1�k�d"�E��b�D��m��K����vO/��gk�\��1O��\�R�JFop��B8�H��2��c�%�=G)>@s���eSm�=L���S�s���a.�p�
��ky@��ցb���f��YZ�@�ed?�gv�:&�|	~M>�	��df�l=����,¡�LYUχ��r����Э>��o����Al[-~R��{�s��,(#q���r*�H1D=s*M�+qqyZ����ū���(�h�'��}��nOsf��V���b����n�9��TԈ�E�G[�/��Y{9�dw����^_0AY[K�Z@�+&!7�m��jn,�6��q|�t|f�.w>�����ts�F���O~%F�=��C������rל�5�4� ���'p��׶J�FX"[옾�TE�Z��Z���x��m�,a����ʍ�ϓ�I�a���
tV�*�_�)���]O���^D��s��	����u�����q���DG���h��	���~׊�`�!����?��N1H*%Y����{���k��S}5+��6_�LLwS
�˿�d �"��
����:��&~u�2��p\���]�C� u��t��L ٳ�?d��e�{�,����}��A��`{EǇi�ץI{�m��x��m���'�WE�/�������Y@[�BB&��읫U5�����cz��"F���O)>`sq�T��m���~K_{<���RF����B��K��>����Ø= �'�����\�,;�C��أI�R��WS"�Zj�1���K�}����_�~�ό��6!ű�����
�����b�T���l����g��nL��8��T�y�ٕBt�����I1��a�6]�\�nf��s��Ā2����25��ܛ~����9'����h��%�e�I���!r���1oB�8iTH����_@�&�E������_�M�����a��ݮ�8h���:�B���x�ao�飂�{�we�͜�2J�2����eo�o��i�)���@���!�J�ڬ�V���I���&���E�S�?ssɁ_�����j݇X%�CR����0��KJ�yd6�a�xi)pi���*��{$�8�$9��"���;��z�ݏ\ޓ�FN�X��T��-��O: �9��>(�����տ]�ο%j���V|�d�;%ސ w��u&We��ה�"�#v���F���:��@��i�p�2�|�9NY� n�G����+k�~H����tVz^o�j�{�u7��������g��q?������?��q:���'}c�����=���h_f>���o}(�}!q�	Y+��i�2���~ �;ɏ81�Z�����q���j�����G)��h3���i����L��s�2�ȳ��=�'O�ú�*���.������!n�=uƩW�R�P�4t��'pL���p�2�;�s~V�W��w�R�MB�b��Ƥ�QYq�R�{0�x�ɧ�J���qq܋P(����n��:�ν�#Q56�@_�NO;=�- �K#�e�7\���k�}�(�~��3T����� �U1E�`�D��r�t��*U�$!j����N���dF�.��(���F�z��A�����U��׵�K���*�i��^����vr�D�t,i����G�п��@Ӷ����6��y��4ÿ~�6
���V��l2��Q�9�7�ʭE�5�R--��r`ش��87�D2+drt��Ye�����a��L֢����Y�۵j D� 8���2|�OnwS���k��u8��C}]��ؔE:y��d��B��F<�D,������ّ�44���o�`=�mjDѴNaǶ�gi�=h�����M.�Ʌ�Auy������`��̕>�*Y��U6���`�AZ �>�\ϝ�(=T�'#O-���4R�S��d��z��Nة��� XLe�W(�T1�|A"��؂��)Vh�8KIXap�W^0u��J1�YkгY,`����޴�T`ؒ7E�]�^�H��z@ ��柛��8�_W]>__抉�prY�^��|7�ai�̋vwO5�N^2�LQ|�	%����>3q.�!�7�[����,���v~NS�Z�q�d6�p������&9%����i�����|#!M�����?Q���R5�,iVX�8J��kF2߮�Ɉ����!��S��Č���E��ܐ�*ctȲ�*ѹ�	�]�o��%M$�\����~9���~K	�8�+�#����Z���z���[�Zt�$��K�|ď|�ѐ�d�┙��dS�Ci@i<��)/�V��ԔN�@�.k�V���兄���j�w$��-)�߮(�:���.��O�}���i7p�I��4�.)R>}��m� �tb�a���E�V�38_nl�P�D�CybO�Y74�F�I��<X'9�0K��v�U� ��+�� �`�.�E��Ҧh�@�4[�i��`0ڦ��l�l!����tc}W¿UI�S�&1e"<6_Oc4xY���X� Gs?'Y�CP��K����gs�ڈ9�2] cr��Yz�T�	k6,�0'zS�ʉM�ͱyfP=�ɶ?3�&�w��,���[��VL��l����Ё��`�,�q�I=�|��U�� ��wt��4���%/r�S�&w��@�ݍG����1-�����8h���ho�\�DHe�d�T�`k�iG9���;��zl�Bs�f �$�hB����%З;�ٞ1�sV��/@Iڝ��A�����}�x�pN�;:�)��2�uP� R/{X���F�����ܩ�;�f�S�w�Pv�G��.7��W���
M��*��Uًn���N"�Ƌ'KՃɢ��q��h�.Z�}��@x%7d�Ǌ5
�e��(�%X��ᔍo�~ �#�3i�V�빔��M�_�@�3ȇ�D[^c,����b!d
ޒ.�PH\J�n�����܉]��=Ϋ��7�����5g�e��}j��t��ʪ��9��G,�$��,+|ax�t�g$1nU��e��[�g_������$��=��W�y�Z�!J����#�C,UŷS�ގE�����6��C���&�1�cwlO���L;s��M$�O��m��y����X�
65.ф�Sn |5�_��?a���k�E�r�LE+<�v���Z�~�۩���%A􍪆Zh�����M�n0��]��'mH��"�A`Î���9ʐ�K��D�R5ѳs�c� �H�QY�d�E��Wsdf7���L%0[�����@�"���A=w��c��ua�]���₿�	�]Iأv�狓�0Ew�Q�dI��x7�ZY>q���;����[J���-����P��!��V>.c��j��[]����NQniv��V��_6Yp��V�����Zf��E���=�0�B�o*ώ9N.f,�hh"�t=i��mv#x	gk,١ZQ�@G�H���d�ܖb<���k�-4�a�nR��:P�<1�����	����ݵ]��ӽ�qZ1eJz��4{�a�}��|���<���-Z��N�|�Ǝ�5ԙ��ɞ�5'12�����w^�w��R�Q�����ʧ��[���˻_��o&��6 ��5N�s`��n�$�YtK��i�s��++`Zy��N�k��c�ۂ��Y�X��=�o+Yau�#���#�[�ڧr+:ү�����R\$7�̗KY<C;1n6��+�5�D��?z�.�]�*����11_�����~�mQv/�KGei}b�%2^;B�l��y��!$h��X/�W�3��cn� ��=N�w���k��Z���������r=d ��=4~��x��_���s�-I^�Y��H��`@*�|H���h��ȸ/�ҕ������Ȑ�4��	�ʄT�K���ҳ������W�����s���	������+��,��TTD��(=o����2`�L\m_&!<5���7�x�@<8�@�I H�(Ӷ~:������1i���s�	��V7| ���'�k��瑓"w��R4��B���e����@��w/�k՟S�����Q�&��D�@���6C��=)s��/kQ l� �!�lDv�HϬP$�;L�d״Z�43g�I*�+Xc摖v�_�|�[]G�k��4��Ǚ�}�9B�Y������J�u����7~��AP�g��LR�J�������{2Τ�r�4���.A�(3�M�#_u��yq6mjbP#�W�!Ci�&{�����mBq��~���"]T�����
�q6/�/oYm�{����ևg�Z��CH�n�RٮnPi�<�oߕ|g��_�pTI�;z1�6��}�K!������n�p	�y�С�^ dָ�?h/�g��f?�ף%}a�&�F���f�-��E B�z/c8�r��D5���Xd �Dxoo�ƽ��J��6#�elI���s��D��]6�^<��L�������nW�.^��zV5��ip܊��@_����n� ������@�'�>K�D�`��R��m�oM-廓�N�/���]=����-5t�"�\�rWⱩ��0BC??EU�#ϥp����lo풼˞�y��Ç��<�8g>���ՔXEn��M��kru��Bf�4������u�?��V(<��%^�q;Qa^c��8((~ED��>\
S���
0R�B�(�%|����(�܁�i�*�R�N���y$k�����ܚNO������}�:�'�؂]�̒GE@�ǫvk��!壘�v��燑��sY
	_^�"�#�<Q�x�~�1S�Am�/:��B�Z���ۮ�|�^Å�P	d�AI�2S����]7f^��^R2I��P�
$F�uݙ�O���o��Qw%�5E�L_8[g���A����8O
��⫏4uYi���2���P�+�����z��>��^��8����c�1�l���Ǝ2#�UqSNZ���i`d�<�Y�?~����D^>6��a�r�3�b�|{	'ߗ�I0+�ǜ��e���2B��Bξ����Lz�=�摒�#SA>�-`�I� �9��DfFvX���ߊ
����ޭN�L�������# ů�K�?�w��j'�Ձ�}�;��s��|>�m�	�
v���v�rf��>F���PE�GVi:P4�|j�4��to���/']} �∣]ME�E�F;r��o:#uxRG��j'��f'_^�~ǿh���\&)�A:N��c�$�Xd�J/�~/a��B�����^{8@���R߽�qYg�	��9'.ɮhk���Cq���}��U�����4��b��M����)�m��-s��cZj��P!�l������������4�eX�0�}a/��n��萖|����0Г5�`H���4e��rne�`�
M3�s{#=X�`�.�_��
��8z 3�)/*#p���e��e�~E�	QA�4r�B�3�3m|��dn��I|��r�v�$u��q�9�������zqpQ�L��u7����;�`M�X�Z}�Á�D�{�W�ћ~h�p���g#�!.����T�v��р��f���jޡOjLu�q�b+���f^�2�/|j�V0;����k�z����:�m�<(�9"����d!\�Ri�Q� �	�����v���@BR�;�ߊ�q���s��f(��i9\�men�y���0�ޜdLܸ�N΢�M��f��t�,�Q���a|�'a�AHK������5��;��t���3gM=��V�rk�Mf��H�([�u.<9�Ys��T�z���']����ؔ:NLo�j�d����i�B���)����)��A)ALQ<�r^W{L�D�j6@^�`����{r� 2�	"�i	�
�3b{*1X����_]��Y;���.��+Py��c!��6y��vO�z�i�Xc��ΰ�u�-������I0��HW�}=�~ڬ�q�>�(;������/�vϟ:UM�
V�>��V]zlΐ�LE�b=s��<���(�C�Q����@�!H�:�9r�i�� V i�Ŏ�i.�)r�(@��d����d�-U�5�F	W�N����*a�
�B��esS]�\��m� ����B0IJț`���w�Aٴp}��б��:*�pSS:�1�s.d2�GF��ܪ�C���=��6|[��Gy*\�z5d�ٜ'��#3z=�s�v0�����	�p_�<w�ݯ�rs�IլJj��{�M�#-��y�&.�;�E����?Pz�6N�V����N�(��>�47�����L:r��E~���,R��0ͤTdiG��rҺ 9�����ސel�|5��8�� �$�4����ڶ�U���5҄�~��w�dK=P�56�Du�����p&p�| 1(������
�>�ݚa$��J��#"5�69���� /:̆ui��&�?]�����V���U�������,��F���c9��L.���+A/�\�%�f9�T��`���a>C�
i�k��>ÆGGN�ߣ?rH%<�9~γ!n5����K!�*s*��)C�(��~K`Q���i� �^�e�W�婠�W�������u��K[Fl�#ίKġq�j�,�&bl�F�P��26OWIQ�Ĳ���^��zߍ�����R��F3���S� ���,�Grqӱ�pA��o�������rB�>��]�8�>�ē�P�dP��X@�.�Y3%-}�6aA�AJח�2*��rw^�nYp�%*�F��d���fX�{of�$��}(6^�fe���H���x|=��_�㷮(/���2a���N�F@g
P����*GGa������Y�d��KЫ�>i\�)C��'��,)���j=�������TE�ҭ3�\�G;�v���9EZV	+x�g}�8�ׁǢh]U=����B*X	ǑLJ�QPs���K	*�N�Y6Ե�^�~25��4)��އ��O�&�be��~ƀ�C�a�K�� /^p�2�y)��輠F���
���7]�r�{-�u��$�;��U�[��5�C�4�9�6�W�:GrJM�o��}�rI�v�`f���rs>���.j�$��/<�Yշ�S-@�+��T�bo�U �b�jW$��\E�f�4{�?�ch��6��)*p�S�q�����3��M�d9W����Ud�G:R��e������kP�y	*cyL�������W
1��{x7N�+�;���H�zE\����([|�Ym��R���T�zX��d��3bD�����`��K��Fg��Z��L��C���~������ ������o��&���{Q���+�+�V��H�����,h�������cv��t�}-F�m��(��S���}ys#/!����J�!'��ʟD�B'��:�4�	�~�:�1/++X�05Շ��4g�����:�1��\��T6l��O�w�~�.7�B���-W�ɼ5H �
�]P�ϩx=h��$t�0�����2(�	^��H�_2m�o�3��f>�L��.�{T)[�����M�Ğ3��9Ҹ�[�7����-q/�U��MOWU4ɖ��"�rm�F½�&nq����K�<�Hr�Sk�����4�ٖ9`�}^�_��.�!\3v?��gMj�s"�Yz�+�f�����y)~E+/q��\G�m��I^��J�Uk��g����쏂�����ӝ�+��?v;Òň�~�95�P�|��[ǿ�aڤX�3j�+$暈x��%S�pPġ,��&b�ݢ�ǵ���۸Ә��Uퟃ�Pk@�&Lb�o�&赵�Ǉo;�����/����Z{	��w=�)�C<DqPC�~�h2*_Nڞ����0����W���>h� l^����V����I�^Up}���7���-8)�ٰ�C�H��Y֪��~��K8<���M��Rw��^�Jk����4���mX=���~'��a�������k���}���[g�V�E�SaH�E�1t�Qs.���7p�u���@Ol↏��`"jF�,�;�'y��ޖ�NE �A����b��.6�����ob.Ѿh�e�ϥ�"~aQ`�����¸���ը�M1�#�.�1i]#V�˞�u��Z��Ƚ�C������ޤc$4t��>�l�3.=l?��0R�M��:��>��l�ER4���쪹2��2
�V�J]W�?������
4R��Mi�@�.�aDԧU"��J�)���l��_��sJF�khK&<��Ԏs��ry'h.��b�B��U]�#�h���̳w��6�N�7EFo��$���
� �OQ��F�]�8Z#�
��RzR���}W�G*���27gmG7~:ȝ�����m��D���^��t�a���wr�\��E���t�x�� |�H����B`�j����`��G��z�g���I�\F1\l�\�$�@X�4����Ĥ}d�>��G�i���3 @��� ��3���s��(��u�?�3�fT	{����gV4��j�m7��QES�L¨��^�{�s	@�/(��Hh��WyJ�D���}�x&l�}+)ɶ]�*s]ɦv3x�*��mO���4�[T�R��i��F5ؚ������L�3V��-��r�_��1 oU����@G����x%�dc�ZSۙDbY�W�ai10�^j@��S���Tc�;��*���Pq���&�S����e�u���������5��!�����̼wX�(D��é�4��!Q����0����1����|���p~���u�� ����DjT3՟0��i��]��j�p��-�Ù�����aI��Έ�~�Ӹ�Td��;.Ԑ��N�Q����UC��{A��h�mH���QzjM���x^�ؔ~�M�T�TA�a�h"�Vv����	�	70�r-�ps�D��Ls��{0bZ���6��]����cg|l�j�ܤ�Ʉ�-,�Q�.�T~�e��a����И���UU�#�{�b�;��~7�p��c�v�AG�_�P�(�ý�6��5�,�PԪf[�������L�p��2 i�C͓P�`I�3CW
_5�Ƹ�1�g�?�ކ���}e��Ly��3	nK����m���hӑ���E���i|��EQ��<��6(�r�(�ZF���]`������J�^mBa��2R���x� @
�ά��w+�ؚs�J Ŀ=G�/�<Z??����ر�nɬ~��K�d5@�$bYm�[�o��o��9�N.���y�ڕ�1]\��1��
#/N�r��~��DV�d��MI���5��,59�U���ƹ4��*��O�d���_�(�VS�/S�>���V�s9��H�S����Hf?�c������h������?�>������G\���|�Lj� �]��L�Е��,�=�G�a��"A���rhT��]J-��i��
�j��Z�=.4.|�zdk�4��5Z6~z�^~�w�͈-��/��g_�5�7���y�^����~IT���^b(7�xEI��5������Q�i�ûf�+T���i��k,�~`������jM�A� PG���Z�|lv�5W��g���Pptvz+�R̚=e�� �\��᾵Q��H�6�i���Ǧ�Iw�8��T�k9cѮ���g�ܕuEr:i���e=��kzu2�?~zl�b�cO��K����G�l7�>K�Z^\+TpT�⃧�i�M �+$��C���ܜ|;����oV+���Zyf����0��f{���, ���$nz�S���rCA>:(�?o�?q��<��T6��RޚHHd��H����N'�r1)5�vG�:>����{��ʳLqdY�/h�v��`ĕq
�'�� ��V�l��TЈ�q��?(��_��L\�F��ߍ������E��{���u�a���x-Vpw�榏�S�n�M��8��ޔ��u<2(�](����?ӊ��wx+�e�s37V�O3��*w�kk�n���>@���_ �#��^(�B*����G�Z#�I�ɞ��e!�:��9��YN����
Z�p��\v����-��h
5����Ȯ�l��!�u�>��5����CDc�c��⠎3~�i=���g1�
�������$�!:��H�!`��E��8+6f�Am��W�ހ֤ؿG�㼉�$x�qty_�N�Q&4����������S%\�$R��/3' nS}JT�����GJ�Q��vW\a�h�}j��;6S����F�
�շ��A!��~�xY���+瘡;R
�c/y���"���%	X��*kC�Iv�q�rsί����ͣͫ[�i�=4r�������.�^"���mC#��0K?�p�Ȥ�E���ws�X-װ�Yv��]"��&�6��P�p�)���"}�?�r���RUrⳚ�}�Gjf?�4K��s�	��õ��䀾V�v�vł�>�
�4?�
�EUX�T���nzig\�{d	��WB�U��J��XN[�����}A�DG�/Ɨ9�v���U�����2�^����Y;���C3&�=�$S\5�����nrF�C���rV�_4���[��X���sA��(QG�>�[���?m��K��EE�}��T.rO�ݔU�٥�֌%0K3K;	��U�C���/w�uN�do�S$}��t��x�1��)ݐ�nB��F����%L\�<���E��7��:��'��}��Х����2=+���8���I�$K��\����`Ɛ��~�K�<%;��Z�sm�,�7&I��q&
T�/~PL��3�q� �7�H�4����z���ȍlt#����HǤk��~h��z�5�|1�W$��L�L2~�X���U���n�*-&�yչ5���mh�&S����1Z�"?S!-/*��9�K�h*�m�C|!� iN��*/[��/?�g�\Ք8"ힶ0Tp,Vۼ�/��q. �"�;�8%��2��c��6
�sW_�ױ�
�����=�Q=_�ƌ	;�W�V��dyn�fDc�z|���Ә�����!K.��e,��{
�\z"�j*�9�ˆ���m:��EJ=8!�2纟/Y-����y-�&�o�M��i�,�d���+'�9+�����ց|������.�g�ꥤ�C����%NkA�IK���T�Z�J^�������ZG�1,.��(��#t|�H�c6��//�}��n�6(|�u$ �:����r���59����d�H����J#�ځ��]�Ȇ�N(��+]~�?��Ӎ�9<��GC��>Po��SJ�cA�-�5���+S�ؙ���s��N�lK�E�J�ݵ����g�נּ�8���]㽫���!�"�;&Ѧb�5ܥB��\��+/�t��
�za`y�oi�'����;M4�$*�V�qx_V�_������[���%��r2^p��<.أ��N>���_V�[6���%�D������qc��M�H%���(����D��`*(	���b�D3c�A��S��h�~�s��C6�S�n�3�1�N�(��!��e�Ձd�53&�Ԗba��>�[aϥP���O��s���" 3�������S�Z0��}����K��R�<~�#�Z���(H?�+�$�'��s&hl47�k|h��8���T��e��=�>"m{�ݩg�������F��vl��u�脈�/D�z� �Y	���L��asO5����*Ԁ���L=M�g����C%�%���ɡ m�+ikE�R��z�����hg��6U�������=�K$�o��. rȱ](	1E5� &F�ƤTֹے�0b=)�.�f9D��!��¡aTX���1���֦����,B�1;�� vӃ�t͔YՑ�?�a��.�,�i�����zQ���#x�<G�R'A����^��H�����B��w!Wntc6��y�TNЖ�8bg\L;�1V5f@	Q6�4�H��;x��_\:�2#Z�� ��O>�C�Bǲ��_{$"��]8Ě��0A�>q�/��1Uv��T��2D�  ��<*�����6��T>g����bQc�ځ�&��[�td�_C�l�T�*�fY�l��:Tf7̫v�9o�M��y��z�-DI��d[�ϟ����Kb�G�!����	�ݕ��}�����]]��P�]:���r�7œ0�凡S�o��Z8o(UX� �J�<D؄�d�����1C�ݏp�nBH�3���n�����Y�[��m�c	 �o|��vGX����7�-�7lޗ�
p^��/¼7��H c��j�����^ۓ�<5F�U�@<`�Xyz�jh*Q�V�>tN%�l��T���=���X���SRY(z�)�s��]���݄�%"`��0�J�O�EY08g��X��M�\�	��VA[1����#kQ����.(�Л�}OQ��V�X�
N��@�,�T&ً��ܮ��@p�ˇG��+`&�-�W�?��f�S�i7��֮�]Zq�#!#�u���xX*t'F��8�>L���i%�.F�ᲁ�������A�K;T��m��f�Ճ7H�sS������<@Y-��ǼXU������s�
/�˒p�U�����$(2�F��ыt��Z��(��XSڏ�ځ��K� *� ^��
*��ڰ���]ǡ22p���-(@�f.|�%#L&��I(�ο��a��� 0��x�i_Sꓗ�BPmwd�P�(��{M�&��'l�����y�jb�	�0�j�o��@�	-���Gn�Ð-�9�3)ڲ��%[H.�݈1�&��b�|�cwn��I�S�?a�A�*�n�a�[�.߃�$�4Փe���c!��@	q�-��2��ä�垇c�׺����Y:�`����F9�s�؇J��2��-D���:�[�M�i�����B$PwÆ���@t�2v?_?��B��~]�37�t��b�i$S
+��l�R!ǧ���Ei�B�z#��rT���{���Q�>�BF������aņH�Î�4%�!rr��i�=-����� l-PW4��~e��@9����VEx��۴�L˃��lJI�9^^�!�^�r��R��9��J�\(��5��*=8����[o��X�&��E��R�:����G�Bs��f��:`��`U�����L�[Rq@4�A�W�#��a󅳁��јפ�V֋����堶�<=!
Zor��D[�蹿P��2.�%���J��Ņ6�S�	y�9�~h����r7r�"�Q���iQ�Ff��E�|��q��L�r`U��K��{@)�+��!��[X�l�6����w���4�ˠT��Gv���ߋ�E��U]/臲���
�K��W!z?�|.`&R����'�[�9�gB��|_T�L�2�ۓb t�1Z0�Gp���h7Q�,��]բ]�%�\�=[���/�(Yf��e��t#�bWf~� Q�g�2;���؁wB���1y�leQ?��N0RP!A���KC���R��Y'v�9�mԓg�\��A6 3cn�����O)׍enp�v�Ѝ��!��w�':;�rԕ�Co����@��>��5ܞJۆ��}�O�Iۆ������*�]!ו�[M��LR��<E�k�55�}E�����r���Y*��R;�O����L���C\U�B10���{U�i�p����2\\�YZ�[?��]�;ɠv+�/�8$�+��j{�Ew��J���q���'aB���dIӭ�Oև�N�bck�8���(���h��2������c��T|� ���s�2��K�C�Ifl� f��z�/C�(ԼＵ�e+��ݏ҅��)t����8q��r$���~����;c�o4D؛�xo�b��Q:Z~?l�e�ĔK0�y�a����g!'����$��22�n��)�0��p	� ��/�d������vɉ�����.�y��(�L��ȗ;k�ž�`���5z\�9ܚ��!��%�P�uc�]b�)�n�~��q��f�{BO	e�ۮ��=�P�j(pqO��4x�3W��ʾ��t��I,xM\�j��b�E5���OcaN��t���a_�p�/�����pgh;a�y3�~���v�f��Ǧ��&����2�p�^<��׆��闲M@���e�W0��ƕ~��,^PJ����N���ڴ5b���D�<V�E_GĐ�dV�eNq*�a��Q-���&��F|+˅,M�;�w�����/Jz{E�uLyo)8���î}	1�97��7o���F{Fx[�rL=�|"��m����=��)��bk��m3�T���w@#:���ɿ4`�xcﴴ,K�<8u� ���;U�u�6�5����_!1����Y�r�Ԉ8�g�m^e>�72㮕�꼶�]�R��mҝ�u����X�A|�4�]��'C|Q�m�Jsl]K�])����cp8;g~߶H:P�G0*P�]��Ak��/=����X��3�q�Ͻf�}wF��,��#�lh�!�݊� 5S`�K���F�>��c���������5�x ���:��\S�[%�:��n��8���u�=`����yv�8b��PT���`�DB��y�<�Dhq[����Y�e�A�:��ݥ
��$7]��� y�3�cPO9a#����y�t�mZ�b��Twv�=眚`Qj���<HP8��m�N�箙��eD��枤eM6��1jÜ��Tnw����r"��]!�5wglw�r�>BJ�iTD&�x���~�-���������d6a���J�5�.C�fNI���k�W"��)u��BĪr\��{K�.E�j����ء�N?mK�X���7>�;�fa1��'œ� �H#�*9�o�����!s��з���:sg��k� �t��F]�/X��%����V>y��t����ɥ��bk<�o����@x�3�vݰ�+�E �q�r���U���	�*���L�`��?�z���c�:�Pٟ[�T.n�t���5t�� j�Yͬ�O꼎�!ٳ�a���*y�*�-A�+�	k˵�c�%nӡJ�4W2
��e�?��@�J*��|\/�9ޡe2�E/[~6&�����N�����`�,-�y/^L�,�~�1MI~O������Ҧ'����d�ng ���n3vN=Z��1xЧUv�8а�q~c�il�9�Mˈ�c�S�Nf4w�<�\���V�N߳�9EP�"�fRI�����c`�V�򤊏�c���2j~�)*?��Sh\�����$ǉ?M9b�y>c%�.>W�|�(g<m/�(�>�nP-��d�v�`?�� J6��	��q���5u�K_ン$�?��jM_>S�Q�H��^�� 8�!�4Ѐ�~�	G��R&�ŉ�4}�7=�^��Tn
�Fd0+>����w�Ԣ9�mT���k�V��ֺY1L�~U�C^�a�\�ь�w�ч�QE0�E��1��Q�ˎ�y�� ���B-`0��Qji��S�p	��+r�G����qyw/
t�ҟ�n{ΡvC�S�~�w0�f�4�r:��[��B,�{��N.P�86h�X�}��z����'�2��)nK>z�x�p�f��{��������1qTԵʍ�ShY�gc�hL��<�E�~�N<Ȁ'!hT�d�6���% �( rPfVi٘j��i��P�%dSfZ�M
��H��Χ�	p���߄�r��N(��p��T���F�76¸˧B�tG��8�X�eeY �+�"������J ko};̷%��oX�d�
��z�$�T�WGs�OǮ �*��X�����֊��w-��v,�PŶ5 >)��/��)�,x�#Aw��{GQA@���R�('�]w:W�Bl$N�r�a�N�0*�b�B|�v�O&��IT�� ��h��&�?��<�6����[��I7�@�jb�ӑP�,�3���f���t��H՗�I{<�S����n �m�G��U���a�O977�zԚ���0��f�2$��oz��U�'O�.8�:��(��W%���G�c��Wk�P��
|�t�DN���!�J7��T��Đ����!�I����J!}�b��snQ��m��1�Ԏ�=�s� ��L�H�3.#KeZDܽr������9���P�i��e��9�v^�M���%��g�
�RK���W,��R{�`��H%�,i���Ϛ��q<Y)`��BRH?='�NN���!,e���8iZAu���#Xk���(�Չܮ����^�v8��L�����]��F۳�����7\?���	a��rtQ�5dl�;=A"&�:J�ցb-"~v^l:�q��*�}f�W���<��{���#����b?�;�0���mґ���M��G�k��
����>�Y�n�*��h;�7���P-�A�.�ԃ�G�E�A����e� G�Gf,�iÝ���3QҲVq� L�>y$1���TF;�ˑa��<�i��X|�۽�����İ."��v�X��)moLa�%�P���	$���P4����� ��g1�d?`�h������rB�F�������n­���U*K<�`	��6;b�B�W�~��8��A���̢)Wt�ۨ|A�q;"�e��Q.��@l=}�d�B�r��r�_�r}�)͢��eM2��o�-ႛ��.�$����k6!j��_��rżc������R<�@i�e��{�M>��C�K�!��@�gB�L�5tg���Z����sK�B��fg
�K��8���v�hR�NQ�Q�5�z��%*j;&*�3��e>~��+H�܅��N�c�% �Mhmg0���f������7Qqo\�FV��C+X碽Q9�G��� ��U3ru��*>J�+o�<�M|�?�in�F+�=��͔<Q�-�8�?c�14pYs{L(&7�;��U�����z������SH5� U(�<������qO��)h��)۷�>3G�j\�4J�m�`�)�y�k��[�a2��ư�@���A��Z�7^��344$	�c�M޿�s��z]s.VMf�Y\�H�.@�@�q��8��LM��|����u+��xѐ���F۹ MH������%9�.d�=!O��ƬX\Y�C8�� ͐}�1j
��7�%Ԣ H�o�u�	.dA�J�f�^�M���U��L���h�̷h���
��7����t�$T�d�)�4��s�����)u����]��n��2�t���'�k��?U���l$�c�Pqc5v����wi:y���H�+�l���<�NNCa�e�2��=�bKǠ2Y�
�:y`G�C��qY
=)�z��L$O�yC�!��X3,%f�Jn6g��}u�f5�aF<#N��,�0=����؜�N,΅h�����AΌB1{Zʭ@*>��������OWX�K:��H�W���D ~��ֿ����4�-����_ؤΦ1�O��B���������?�+b�b*����x`a�iI���#vԨ��a��_�**��Gz��A�� a�N�w�t߸JݠM�Z��(;��6*�6��aޏ��4Tqf�����iY�L�uj0�8W-z3������9Yڢ�Y��e��>*W0�'"d��9��FZ֓bBkIA�-x��<Cf=��hņ�����9�	��n�Q'
�\�,����V� �E�oa�cR�,2��J!�onk�4��S�>�}���$����2��8��rK�6�%"B�(��`�������ԉ��K5�.f�3D*x��b��Om�:
�b��淁�wN��]�/�_3DR[�b�ý�]�Eh_�⽺�������j��&��:��d��p��6kЅ�¡��d�6K��$��<�K����D�2�`�-{�a�ShIp�L9ެٯ�][��7>�pNSČV\���:�39N�`K�th�$�l�#�U�����I\�؃�+�5&A�z��rs�\�[~w�OA�A�}�c6!x�>�`]]���6���rrU�1��`5��f��ώ&ڍq�a[�oQz��2��k��Z����Dfd9f3LTCT�f��p�·�.���J;��IX8a���'�"�Es�}�D���ÑU� ��?�ܺ�qn�Я#�޷t��լ� �oBFX10d �u��Eh��O���wcS2[?UKx�����	tX3����,3^�p����?�nJU� �kLD:~��Į�
~� �tQ�I	F�id�}(X�F�x�Y��}lkD���]*mIe?E�p�@��u�ĉ�Xͣmb(��Q3��$�=�����y���f�y�6��ُ̂=�b$�M��˼���0���L�Iᗸ���94m����B͟�H��M8%-���V�@+��� B#W�˿q�_t���G@s�	���(zp��X�p�+�	������P��[�Y�mO�g-�U�貕��VU�\ER�@I����I���*�v��SO�w;��D�h���Ŕ`I�s�\;1|W�ƈ���o�����7��˔+���&!�V~1 .M�e�Z'.ד ]אH*i�K�����Ԑ�%`�����Y�߷ס�bؙN!b�>5UX2>c�ƣU���榩�>En���m,�%��F����+:ϫy㵶��c*̖�Za%
opZ.΃�&�r���[! ]�R�����R.�'���lk��/+���h�1��̄��	����^�|=���<�S��/u��Cv�'����(~Z�uUS��l��0`[6ʋ ��;����4�)�(�?Ӻ+_e�&�o� &��g�<��<ç"S���Hq�Ys�݋��.e7�4��2��^��;+��燶7+�����8ʗ�=�a�z�cM>L=�ҷ;�ી�=�z>��X*#vĨ���M�	ˌBƅ;��͸������A <�?��mbZ��N=?��ԍׂ�͹3ϋ3Ț��m�D�A���k��u.�*4Q|J�4�������FV	?Z��r���M��q�o��a�؄X��~��9�C��c�Gjz���6���ĺ��;[�{�H�B�,9sxƯ5>̛�R�<w)�0k��si��#��z���t��qD�o��%�*�N��������̕"�?H��a����s;KxˉQʆ��\�q(���@�_��>ެ�P{�����/�݂g�@M��S��`�&lWV��5x��tuީ@�I8R'ZsW�L��r�k��i(�qX,!	�~ҮO������ ��#G�����*q���B�b�O��x��q�:�|�aԵ��A��U�KI^�1�3JV�])�,¯B;tf�I�y#|bL��5�ky�=����� ,�|(�d��X\k�������)���g/������Ξ{��V*�����C#����Ѯ}mj��
���<s�ɧh�3rNg���;7�Q
B��BW֩2�ʋ��&����W�d6�GW]3���|�f�0J�/�-pï��aw>c��X��R�0����M=�a�� ^<���^[1RT�cd�'s��-s�����:]TF���t# ��3f�-�17$���>��T7s���w��rU;Ѫ��%z��o/�(F�9��r�6,c i�h��W�*0�����4��M?���0 �H�W`���.�t$���4�FLH����La�q�-K�a���ٛ�7;#��B���c�(?g�39?���L7�j9�85�kq��͞U�&]�&���+�X[,6W�BB�ߧl�]��؜^�Bj��5�r���V��K�|
�оˮ��E��><%.ݧ�]� �0j��"��a鄈�g�A��R�J���3W�þ	���0����f�J�pF�`d�-O����vM�JbxQ��ύ�:���MA�ɉ�-Jt~+�� �'�j�B�o|:g�+>��n@��6�(�/��
e}���KN�[�v��\ų[��i�a,�6_?����&��Q#�Z�~��R���$V5�a��AL�{$i fM�T���F@�b~�:�-#���'�W+���w(��
;�7�U�c��c���df^~vƣ�J���(a�[�RJ;J	�G^1z榀{�2d�
��oN�1�CfS+C�ƃ^35���-fι̌�܅�3�QmqQ����I�i����a���h���>��[��+�ݤ��%(@�J�	�R�5v����꜈�]��~�{ǆ?��+��1�����l�whk���<�f��{�RM���1
�v���)������$�S�M��n�-4���
��RH̩β�c�!��o�~0P�����F�3%�V.ʇ�2��Tj3&Y+JB^�F��l��*2�&�}���Nذ\�'��Q܂K���}S��sL���*rGԢD/�M�>������˲=^:�"��"֖�fy���Z��_ȴ_�����(���B>C�}���½�d���̘�R��ψ&����nB ���Ё�
/�mG��ޏ�FD�����<pSfJe�?�_0O`� ����YrP;#A� ʞzS">n�=_��p?�"
���������!|>�V���,��[ȩ)�h�y�`�aď��A�V�/�=��Jub������s���9-%��;;%\&��a���~;�Y�u�D�"���5�����\da[xvL�����h�wu�ܐ�p��T�_3�υ2`�tM��7�~�n��V"�B��R���l�~��J
n�:��0���󐝀kA�'��I)�T+������'��ve/<��'Yɶ�"=_w����V�AS�=�@J3HDrv��0�x�Ⲧ�-&� ��[�
ſƿ��%x���������t C�&@]��;�p*�ީJu�;�I6����p����_A�V_=]�Ĳ�Y`��x�u�hSU1�ݨQ�-���n�T���ǼhI�*�e�ahO�mA|}MQ����1�4���.7t<Bҹ?���#���k�xA�JXZZ	��Sp�e�R���qV����t��t�<�#Q�w�|�zqIb젢_u���I�a�`�(��B�at�&}���0Y�I��p�@��V����N�nT<~^TI�lQ�LO����N�:(#p��J0e,�����s1Fro4p2G;B63��]R1���#��mkX�d�����j�	�h&t�("�ҠF�>{T�7��ʷeԭ�	�i�ut�rq���;��sӞ��q@�ԫ7K���|�Z�Eu/���(�aRn��A��)��-G�{��}r
^?�Q�[����F�9���^���G���v��3�0�`�� ���?W��)���1_�cT3��G`O2�QoR�'!�1�������e�0��N��k���wB�]���d����L���J����H!�&�#$�}P�3��MK	{��?����>�4�Z�����h]��إ�j�{\2[���Rڑ��AwF��%r� 
5�F��rV�wu��X�m
C�һ:$8��/q��dW&���(��[j��v��-,ΐ4���|������R *dRޥ�Z_��q�������J�H�2�lE���f�iZY��@���q���-_PQ��fQxi�$ݽ��?�$͸�]8��q&�î����^F��)RvY�N���r%�V��,yh.|
z�%Ӿ`Bv|��7��RگZn����tb�^��-�}�&��|�q�V�CPz7�]�%Z�(.��A�������3q1u�E�6��s����B��l�8;^T�(n�/7$r�^)���;�Uuc�tM�&�@z���#CjR,7�������1�\d.{p;B��_�W�������b�G#W��>�>6?�
ҺG?��ѕ��f�;'#��bB�{���致t_Y�HVÎ,�;�a��{��~������˯��q9�q����� ��wb�������CP�Wsp2�J���{&3�	[�8�����c�|���A��²]q���'2K���5���tN�
�L{������v �!P���4��X�m��s�F��0�:��c��g�6:�6���u�2[�a����L�67	э�lůu�ܧ�~����L}��c�A� o��y%���g�=e����5�[�'E�N��o�7O]d����9-}.�� �o�L�5v�󮴒a�쨕<�G_d�n���G��F]��@M@d�CU=�M�!HLN��B|��*9�������+�UE�������b3�meI��'�$}lMјaC2���@��L��4}�<���g����h��<j#�9,r��=,�\*��Y؛�O�m��	G�,�O� !���3U[m�[FS���C�m:k&V��b���ƶ��U.]n>"��٩�`�?�"}kWƁ�[�F�K�%�T1�-����J��~�W��)�^�iU�{�.��q��,����V���~� �E�뽱�ǭO�����W���٦�i2�@k���	�J0���l<ͨ�� |s����Fֽ���~x���.~����lG�����@/�Q�Uލ�]�6'�@dn�Fmɢ�7n�#,Z��jF�=��h�0/춯|V���%�q��s7b���q ��y����G��2�r����h4�Gn�Qc�K����>����R&�-�v�߅|��(Ѝdg�c��&G[})
��0z�O�����JuX7;��e�a�3�ou�� �xud���A#�6�e�ͷ+&��G-��%	�@c�(TF�~�'��ǻ�8*�Mk�x���m��
ik��x�������|��H�HI|S�����p]�N>I�x��y�	� ��ѮSM�5~ �jx�C{z��0C9_�օ8�\�jJ�~U�=�m���@'5K�F��ᵄ:��;�bI�P8=pD̘ۙ��-d�	[�c���o��`��jJaCQ'�p�,t����p�1�����Y6��$��tb�������=7����3��׾W�G�0�IED�A<�
M�n}�L����hN"[�^�k��&��u ~���]t���T��d�0���w��m��`�Q�! �8�[�x�H���'�y�8�^k�K<��?��x��6��a.������u�=,O����1'�*3�J|���p���Dl""BS�V�cy��d=�K`�ݭ�?�t���m[0E!���`��,\��`��"C1ب�K�E��M��3�Q���X��@�i�F7��W>Vuç��F�#���'��nn>�:�U����XH}f��R�&�j8e��2�}G4}�)���O�H������H�O֩���Ͽ�}���]�7�<3�b
__�}�Giz�Y�Ӗ��5?6�:a)|ßw"'�s�3�VQxQ�/�����*3���#���>��杕�?3 ���=�-�D�z?�ԧ��Q���t&���K�IA�D"�d\W��2X|#f��~>�,�\�*]��7Mik���IKM�)&B<�*0a�yS�S�k���4���jKAgj���'j��`��mN�XA�N���������<�V�~`V�<w8_��`Q
�C�#�3��$NuTW�zĉ�h��@n���s L�[�������V"�-�b��"!����q��zy|�.��?��`i+�a	�:/d��OkUj�Ilp���%d	|-�w��x�
���K(CF�:*��l�P3���3�ND}\���k9!S�|�N�B8�;�k�="_�1�+>̐���� �|f�M�r%�$M/a�v	��퇡s�. al�6�}"�[^�`����k7t�^uJ����Y��,y�疍"��L`��U�0��9�a�L����B���Jy�,\�V֍��4`�B��� ){��Im��;��=�0U��;JW���2ZvyK�v����5.�J���M9"Z�����PoI��M)�X�$-U��F�� �+u�K��ag�[H0E#+k������BS&:��&Q�3����H�\1��я/�6��.e����k�qՁ���JΔT�]���ޏ��� �+M���vS�V��+#V����e�Š��Ǚ�x�R�@݃F�ʹSX�?Q�7��T�ٷ�����uj��`�2�o�)�i<E�U^��3��]� �\������(k��� ��wp���8��.��-�\Z^w_8�"b��e̊�I^������� ��qz�6 ��x��xYVE����`F�c.}����.L����S�x��-4��	E�(ޚ7D��+��0$Q���I�1T�/�Ar�L�U��+��t�V9���&U0���Bǫ^�3b�b�B}�W=Bc��f���$���|���a#b-�>�̤=]�"q�ocm�ץՊ(R4��_�oɅ���FQw������zĭI=��RX��r���t�eP��wc}d��?;�b���.���r}�*�����b �xؔѳA������8��M�n�~��Qҏ�g̄dG����E����ݚ9�A��Gw{�|��[J|�B�BiI��#= M�k~�>�Z��v\��k�}i�ѭ̾fO� �C�]2���n��A���D{k��\5Yã��?�9g^�m`#�dY�1�Z���wpu=-͗?W�VU��//T6f��	@���}R�(����	���w����3�>m���m��7�QiI�D5�1��y����7	�'3﨧�S�TU@���J]�XXL�2+S�P��1�R���6�f�G_�C3���@������$,����)�_4���%��Z�X(`mPu�'n��R�d�6��6�z6��Zq=������)�.���c��-J��x��p�t�\�����a���|3x�J�0&d��0����o�f��ݽ몣���%C�A@8�2ve�/��?n{�����?-�������V��s��iC7㾥^���˞H��9����(����I��6��/3��)P�3r!����\��*�5�IJ��𫗐W�]��0���K ;�`<��ܙ�.]LJ�Ph[�0gɶ^��+
��p��HF�'S����x��>)s\oΆ�
����8�����4X i!����~�#�>�M�E�d�B����*�MEA&F�!����	�pO� �I������hpLO���D�ᕠ�7�~y�<k%`��c� ��U�V�E����O�EV�dZ�ߞ���*N:3q���UnJw��]�1��c��Z�����G�����i��4S�y�����>	�c�������#�t�w���B)��m-c��S*���}lK<��;4=��?�VCm�sh��+��(Q���C�]��� �q.+�ꛧk�Rr!�ͳvy:�T��_Y������9Q ܱ��L���G��,��vf+��0�ג��u�L��d�x��k+��L�|	40��j�NMx�A!��%�����t�!�Վ���1���5�Kch�$���>n�H��p{س+p�tUb�ZT|���]v�BrU'��G\TXi�m$�1�d
�G=��MG�"!Va���;�P���A�m��o�>�m*A_��FwC�a�?�sD����������x�m�p���iMc�"<��x�\B5-NǵQ� ?H>���(ʳ�`` ��\���+�.h���c	n���G-χ�fBH�JTn�. ���@8M�\���4�[)V�4�����Ԅ��媓����z�S �BĻ�L�#�;7p�;��#�k�,Z�W����c+L��������D��Ҫ�[M�d�qQ�	�*Ҽ,�eߴו9���j��jZf �?�[�ĸ.:��}A��!��-�2W��$�g��J��el'Ƞ@��4�uObh��!�o�X�>������f<�8^�04B#�����ZV����N����VL�nވ�ڊ�R �v9���j(��u	gؤ+�I�>�wCv�-�M��K�o���1&�e>�6��(���!Af�n��:ꓲ[hИ���1�e�X�ݰfg�{	��l��.F*"��+���� ��r����R���B�AU;��vm��Ĥ&��YW���AYl��62ʆšm��$	T<��i^�k]��<l���-�-y �qu����T��S�~nZZ�4�%Jf�_�>�6�5��u��աp��w �c1X�x���W(�{�U�{A4q^q��(��es\ 5���5a:D��č��IZUxA��Rv�-M�rƽ�=C��B��lnV	�H�>r���0���a�&_��#1�!OoU7��'2���p�>+���9j��7�����~>���C��WW~>I�Q�rWy��܇B�b�"_����Jx%F���onn]ݏ���Ϛl�c!h��Y	�)�N_�9l�\9����#����k�
��#�'�!��jP�x�SkBe��5��PRP��(e3�'r.��1V�d��c,�c�RX���8��/�vDm�I|' naY7���Rsv���B;{ç��+dpЃ�M����"Z�V#e�V�d�����~���O���J[��%�U���#�ʙ����y��[��� ���3:�f������v��t��)�$E������1�6�~}ӯ�����` G�=/0-l\��x�h
)��'D���x�,�-)�w[�D�^��qG�R��>AT���7�>4*��tDC�R��}}����ºUE�>�N�xLA���Nxp�K.�
���<o'{��f��ݯ���}?��(�ҹ���{*=������+1�.F�~�4��e���=���J�Tl�D�=3*�%��E��и����\�B��}�xlX�z{Ц�0��*b��ߓa�<���91i�B�/�oҗك��g��|�Ҿ�Յ/�8[�һ~�%�i]Z��/���#�Y�k ��M���?:/t�D!Uv#Wa��?3�ˀ��$/5Z|���B��¾Iϼ�Ol�����T�Kj�|U@�&K�Q�_ҙ��y�X>d��؞q���oo�sK�1&��ψ[@5�0R������8�cq��,�#�W���Ҷ�xy��ߣ�(g�T7��� ��
Pʸa��V���C�R��MiSb�j0���w���⾐M{K��0_���D�6�?$��P��,��GDq�I��bόR�j�2ǠU��zD�y8S]*{S�?�XV�v�;̀��{)h�Q�t[��� �1&�J#�L����ke:��b��8��	��
lMᜋ�T���^NB#^|>�ܩ����O�j�`�`�[!�[A�A�u���Mx׃�y�p ���
�b�߲�G�ĽA*�s=���'�X��Z�qڨ�+������CN{�@�I?M1� ��y۰y?�E���B��H�m(�0u��_��?�����r���a�f�و��H�3FA�������#�u��P\�Ff��5xyhN��6 ��f��s�&��U!C�2S{@�./EH��t��M4*�k��ʽ<<=��B;TX���/��xų�V�A:�����̾n�	��/OS	�:�8�IP���s�0˦�㨻}��,���^+�P�TB5������\=�c��s�����mB��8]=h�w��6a��;Gz��Q{�����M���(j�nG�$�	Q�Z��l�k�J�Y��=%�%��D�l�@�p�Ȟ7�_d�)�P[��7ꢧT�&)W�X��-2���CS�P���B�`UJ��5u��n�O\Q˙��"������^gP�����3w*a'e�Ț]���#���#",)��e各[�TE0��G*� mj�랮A!��g�	(����y��s�P��S��~��o����Z,���)��&~#�}+an�gB�z��j�}��*��<��.
p֘Xg|��ل�Ys8RD�tWU�n�m%Pg���`Y��;d[�ѣ����`���)C���K �큇��8�Ӟ�\f`�G�y�,�j$ѩ�Rt��AD~?V�|S�N��8�x)����Z�pi���d���hE�[��s��/�z��O~���"�(�ǰ��{���Z^�JwH�%���<��UZP�m�mZ�R$(�@Ʋ�nz^g�b7���Mw��ӝ��Ss,�tH7͢ Sr}��\��*M	�Kcm��}�\nQ��7O*@W��ZV���,�Ϗy	���[��pg���F����t���h��_c�������d�V���ռ(��9d���\�����I߅H-lt��5'�u��+�=��hRe@�uf�쐽�S8��Ĭ��{��LK���,`����I��";��3nN3
3h����>���Z�·�]��[�5��6iQ�f6C��pifD1+��P�n-=�l�Jt>��O�+����Rq�2��Y�<:�]w? �V)9����?��f�<!r����IY�c��R�S��ʌ����?�JF�сʮ	;y̒��O�a�բ�-HK�jֆ8��J���X��Щ����]�����\B��e8�*'{�Q���Ol?4�s(J(xLz�@���lJ��140z0��N�V��9���ϯ׮Br�U]�c�n�܍�hr)�ڍK��rhknȻ�gث�]�h\�`G ��:MK�c
�'	ه����a�k}7B��Qӧ�R��%��~��Ű3�#:guD�z/��؀�5Z��u8�6���s<�H�F�&�Nl��;��d�AE2\��sF����y�^�R�����]�;��s�hRe�f�
�S�vr�h���{	m]%�JjD���a�M��G���M_��ѕ�����	y� �^�-��p�+��>�+�����<R_Ѝf�����\<����\�i�^��<�{i0������d*f$��H.li�A��oL�Y^	]�O�q�k���������	��1��zG�33< �I�g�樻ߢ�t��r�~�As����@�^Ę�wF`�ީ=�bl�"Z�DP�>.���VZ�O�IB�tv��8K;�u9F��/*E�b_l��x���\�з|-���`'�	W�կ��r��eq�KT8�00��]Z��İ�v��uX%�>�s���ھ�?F��z�Kʣ�4���Y���Q����(�<�
ð�B��U���,��b9����q�Ip���\٠��i��t�$h�R%�4����"]��E�I�"�/
Y�cw�:W׍\9�e���\MvHB��.��rLz)�;a��_l�]C-� ��kLά��}��F�-�����zso!e���8d��i1eޥ�]ǎl�ʖn�YZ��4�H�ko}e�����̼l��s��]�$-���]�]��_���x6ܝ�2��u��+�Z�!X�XE�?g{��$lk����L���Iؖ�E����<��&T.m ���=;#�RVIT>=0��r��LH�C�/���E
�������ɓ�""��w��93����a���|��c�����;UA��&�Щ��X�p���+3T�؊��O��:D#<�����yX�*�Rm�(P)����WCb7JL 2#��(̝uqR����U �����"�$S\b�̄��b7|�XdR!�t��Y��<{��!nʀ��غ0$�]:o��n�ȶ�?I)�F��	TR�9=x�D⧶}G����ϹGɅP�=Ԥ*Y�تG�)��u�NO�%.�������k���ħ`�oi�}~�u�G۷NƯ�ퟳ��lbfql
+ꫲ;Ҹh;��u�?)�<��)�s�ʳr ��쯴��Gb�����i�`*�RzX�cg"�:����<�^p���to3����O4�:�#㋓�\�ڇ�W�F�L��c<O�M+�����[������%$�v�:�o�.'=\}���>O�c�'��A���[1�2Zf�&)����E�r�o�&��<��N{��������@1)�`�2�'�Bz)ͳ1Rz`n?�L9�$�G��6ەs��g`	�_bW��Q?sG}c�_�T<{M�$����	ڍsepe����f�R˩�d�"7���g��8Yw��<�;���Jޡ�s�����k_�Q�-h��L��j�j�{/�������d�yX�z~��X��'~t[�~��E�&��l�g0�咯�� �L�	
G�$�����T> ,��w��q��L;&9ӓ�S����6��{��A�d���q�I�2{�^�)C��o����`����������,I�77_U�z;��V�bk�g�5Ԭ����SX�$��s�O-�e-ϥ��E�Lw�vB�\޻|�j��mx��&4m�5��לV.5��-u��1@N�c��Q�a�	
�-�M�� ��4�J�1ӂI@�6�����ey�Y�]!ʿ����[�hX��	E�*�c���$�C:�����.��E@�����`K��~�� �x����OK��_o�v]N����5��2����O��v�9~�j�⦖K�O,�mb��1�Y��w���^�ؗ|[4<C;vj~۽~�P��ӟ;�/]�Ԙ;���~�u.Aܛ��!��������L �{X����0�%���x/���T�s$y(��E �y���&N��Ҕ*����ts�VW|9$�M/Z)����L����p]���G�G��V�$tO|�a��\�F=���&qk��mn���	cOZ��H(63vgRv�WMB\i7��}��ċ+-�Y#��1����߶�̦�� �aM`9
R7p�w�������u��?�����Q��I\��5yb_�qN��[��T{��z�©����[�����I����u��Ĵ K�����'Pf%��$W˚E��>b���o2_( �p! 
�זh�dG����iu�w��	����MB"��Z#�V:�~N���X1x �	u�E`�Z��[9(ύ�;m��f�ŀ����:vk�F�L��F��*=�U����􉕸[��p����(�zp�,:�}����,^��>(��� ?�Vȡ���Db�`[\�^1����fs+c�l���)�E�!w�=�7�%�:�e�ͼ�Y_s:�xZ�~������X��X��l�� ������ �5A�)��"j(!�m� H���9W�p��J�L�?6v�mM�6�m��5�24I�]�d� �����������hW�ϭ���L)�	�q�c�%K�bCuu��Q8�n)E���{��^-l� ���E��9�<g�(�Aĺ�1ݨ4�H�w6��D& 	'��v��Gh�� �͒���T�e{�|ܮ�P� #s��Ln�P�����6xO�9�5��B5�K�;���gt3�e�`8��喪|���b�䟁���h�x���2��d��	m�\j�=V�Y0H��1��`�-��&�IO��4�^i<U���37�"|٬��s��ܒ0�~�!����d�=�=�}A_!����0����@��kf�S7͠�g���_?<+��@�٪;:`xu&�Һ�����K�q�'�O-#?]f!�3� <|r DR5���� �x�?e�:��z�p�҅(���~�v�J�;��@���+ğ��8���A����M?��H�Z��$ [WZ뤛g��>�"�F�L�G�i�)�ZE�;΃� �KM �i���KX��4;�s}Jy����ôWY�l�T�����ۧ
�{�R�&Q�N=��eNDs.5��QP,�*������sJu�nP��K������:;�ih�Ha�iB�u#qK�jq�l']8w�s%�{o5��7�(��:P�@��ƀ��)� H?(I8���ݶ8{G�l��Z�=��3�� ��kN~<�n��lRq�cg'n��ca���G#Y+�`��c+F����ս�|v�|�xTza�w�Ia�Qf,��P�xň��a�t'ӈ�L`��˝�%P��������Z-�k��ok	��m�-K��ϙf6�{��HEy%juă3��Cڢd`5�g�}ٷ�={�Ũ�V�H]B=$�
	W|�ߙ��^���b�d��0�/�h�	9�"g�af�<��7�H��_����Ν6�!r�%.;�~��`���`$��F"E ~��j���wz�D�	�%�:'>�[�k� s�dSy
J���x]�kk�H��8�P@�����O��̺���8$B��ol�a�AY�7��yy�8�g�v�9�_�!�	[�f�35gyH�p�5��*�hȀ��(�+U����)�M�BR0^��y�v��01X�ˁ��՚��yz�7H|�R�%�34Uߞ�=�C�%mI��m
��bq�������^� \���B�PC��;�ɼ|B��� _�I7��-=�`�K5"!�M�����S�7|�DZ���V:C��J�J�j���q�����k�˰-e�̚OR?��˛n��xb������!oi�V��� �J"`u��f��Pyb�5�?��@��b�C�aK,����@�9K4W"�hy��g��՜P�����F^���(e�&��6B�j���t�����˗���p�V�ڿ�E��V04����˙��Q[����̠1�t��]nX�T��щ�\�tt1w�Z��L$�H���j	G^D3L�Iig��~����r?�O$�Xˇm�Is�ogИMօ(�Z5`�&�_�ҕ��r��=�n�n��W�6�CS��u����ۺ"@�&[�F-:�,Ik�U��)x�3z��K���q�!�5rW!��$���첁1���	՗��p�RĀ|�y�=����<{��DTc�1O�)w���*"Z�1?��i����0}E\p}u�[y�Y)~C�!�\�(ٯr���5	^���;Bk����f%nTR.�v�����Η��F���C)2mkſ��z@"��dA����/�:��V��YMC�C^T_�j�"���dx/RK2���;Ƈ!C&�ޚ)=�)Y���,U��B�l�xzp��Ǟ��.�k�ɾF�)ׇ���P��dEZ'��gLޕV1�9�� ��0����IKt�^s�"W����o4��Ec!r�
���r��2^w��v7�Fo�|���q'�����4�.붞��z��C1�ȓ���xkR�4�JOz0���`z���?���_ �"0�U�C�sZ1|Pp=&�{4U?�啚�@@K��fx�܈��0<C���Qϻ �h	���e-/ݥ�y{ ��d�;��;s,��٫�ڏ��Lw���w��زׇ��L��?��
��v�O�)(>fˉ���z�K��4m�Q�Y�҈�u�|���	�ة���(�<_4z�LU��l1��Y��m�18S�L�Z˅D#�/�$+�^��Ԁ�<S-��~�&b(�ܐ�?� ��2~�ǤA� �e?���*��R� �IH����	gOKڥdQ�+����m�S]�g4�T�,5q��A0r��A
��u-'������P������p�%ڼw_��ϲ��GǕ���P(S��c$^��/�z�8�fqŕP����F�4�D�\�M�j�?��uȗ�X�-��\i'���\�&R�j��ώ�¸aC�Bŏ��$��z������ԔݿX����c�|�]�w�>j�խ����B/��TBSV�3���3�|�)�����j3�W�ߌ#�M~�I�u\�R"h_FĂ���y�F�ޅ5"����V�=�X�o`��k+�!�Վ�q�����=95x��C-:�k�
d���DT� ���R��\S�%�M&(���Ç�_(�D?W}κ�n<����s�L9ۀ�fd��>�����n��j-\a7�#��W��]{E�1Y9���;B0t�7��Z~Cd$m�K��q�b�]S���;���,^pD�~uz��X���Z��*���{C���G}�C��z��q��\��nu����^���F����H�o�x���)؝y)`�ʈ�H��c|�ݾn��i�5���$�Kx�xi��I0���'O>b.iT;��/cŌ,�U�'P�ͪJ��`�������h�r�.����x��=�ZD����Y1H������6��;�+U3z������UYxv�����S�z�01p�z�sF�Ч	 ��sD����I�n� Gs�#;g ���\��n�!��	��'��!���#5ѫ�q������7�����RmsV�.��l�-��>�/����;g���o��`6y�˘F��{�p�4t�ҙ��q?P���i܃3C��}�M�C�A!��W��=�����;�г�R�
k��6�ÓG0�L���f�E�v5/G���Lse.�f3�H��RD��=G�9�أK5�3n��l�lŋR�xjj.H�쏾,��^�4YN��K��!�Y� �
nQ:ڒ4$4��\�V}ȼ�E��G���8�>��N�QVO���{l!��;i>]yH����P�%��4�Z�~m`�~`{[���(X��9R�B��[�De�FaWg�<;�����bZ�0���2�\�����v�uA7��2b΂���JRI7&������N�6�0���3*J,vD��Fz��{5��%;�dܘ��_��	%wJI%V=]�_�TZ�O�t�5�Aנ���t�u-�gB���&�-��i˶@_׃#�hE\y�]�6?t#���*�ab�+'�W�u�љz����Jb^� �;��������͂��.�b+:�Ƞ_�E���c^��)���~��E�d:�1�6hkSW�N1q��[ר�8�?V3���+!�>�$���f�_���˾4曋Bޤ
n�h��N*��y�B;�笛����im���k�@���AIhI�����h��g�y@�4e��|���n \���t
�b��Ay��e��|��W�x1�^Y%���N�
1H���5�\�>}��0ϭ��H6�+-n�[�r��[��G����(��]�����5M'�b0�^!���p|G�ԊM��*��Y��k��GK��<
��=ĤI�5�VdW@|w(�o�, �����^��g��D���K?R5�;dM��Q2H�U��s�)��,�$��y�J����D��E~Ҙ߱ꗻ�PM�aI�Kw�B���RF�Fy�遞�bF�S�^~(И��B���C�Б+�o�i���g5h.��5ү\���lib$o��8/>��&���<����i��E�3A��3()\Շ�;P���6�`]�����A�����(B���Jz�j50��C�/�O/�xl7�fp_���o�u�l�\e�E����UG�Mã���?���<ڶÛR�)�~�h8:S+�T�����������ܫn}ҵд��0�p�:r�t� ����� �?a{J�:rP�׏`�fWf_σ�y�h����X/�{�L���Js�$=��@
��(���8��?)��gҿ�}Ћ���N@Cȋ84�B�k؇�$	����<Y>�QX\R�)\w�����_�n�K��A�kxb�78�Dh\ �Zmc�S�S�'~����=~�I��X&��0@9�A����3����'��jm��csv�Q��=x޵8�d�L�)�q�i��kR!��3������r��f���k=�M0��է�lc7�
�m+��n�v^�f��"@���f�0����	y�Tf��hJ= 9���-/��tds�Rܗ%X��ݔ��mv#�0<�N,�=j�j=UrT�y��2�v_����˽ jB�g�"	��T�(J_�`�G-Zy)dA ��d0Tc��.�W��,S�cF%���JV�_=t�=D�Op��4�m-��/�~�m�s�'H�py��ui�CF�_,���ze��UN���%>���$�_����yFi���,���Vs�?M��Ҕe��r~�w���!.��`Pq�$���r�E��J�9��=8�
��i�x�tg������C����w��F;��[8��P[�+�٬_J���m�����l�C��h��x��c�GU�s�F<���1a������"��2�fk���o��E��?�q1ʖsb�<��R�]���d��Ilqi�`4��r�Vr�s�����W#��=֠�告����~���O�є������P�lO����&�am���_��5��42���d�I��z��ұ�~�����\8[��p�,8
�!oğS-\×�i�e"55�sN9+ o~�B.��"8	3��.���%=j�K^L;P������:=�� ��{���9��|��x�~�FE�����W�5�Viϔ#�O{�д466��d�If��ca6��]*��)��ڃ�g�`s�Z�����]3|�$n��4�c�\�9_�F��_�&;��4�/W*�mۓH8�!�k�*�'�j��b�Q��T�Y@��I��.]H�O�[�Hh�Gc7ޯF��"b;�13p�(Yf#)a5n0�^�x�%�#�/j�y���ݍ.�Z��/�"��7��m�mփa݃�A<�rkd��HsM��BVY����K�,Ilyjm.��3��;�>8���V���B�=�[$�:�[��T5Fk듀Z�iN�����Y������$�\ϰ�Ԕ�{� �#�6���/�c�t�,����if��*��S5Obu���}�ʏڈ�5?VE�蟬��A����+���8�7	��F,/Q�9�6G����y�@�T�������;���=�E���L��}�h&���˞U�Ϣ�3;����\����oR�� {�c��-��H�m$e���3�{ɍ��e��g�Z��A��J+Bq�Q�@�ɞ���Wy�a~i�q�bx�ȕI�BῦE�����p>�)ǅoP�]n��	"�U���B�% �4��T� #Xe��� [�����)"�?$O���[	�s+��k4l$6��݌L{27 �g���0ܮc�����z��m^Ty�}��f]�[���c.ꝊN?~!�h�8�TP�J`�]O��V��O��3��K���d����a��@N #S���߬��(7�ɳ4���w��gݴ���������_��ht�v��lS��3_w�&x	t@�nsm.��� E:���Vw�́l��0�xԂ���6,���}W��:Y^HeV%ݓޔ�Mq+v�%��[����*4w郯C��y^�-#@V�J3�*�����Ѓ_.����B�G�@L�)S߆ � �QbvtD(�ԏ~�K��|R�=���\����@d�Ug����� ��,��@�-̷+x�v�)�Q���|�;s����~:*EK6?m�Uk\p���|ҫ=6�]���i�й��t�y���;W����C�h�`FW��Ύ�uQ�c�~�mex�q�����Z�Ew�@�YЏ��-_����u/�L�w�v \/�%��N���T(�,��>S=[�K�>P*�e;�����lp7�\�7�1w������Ň�o�F��C�)n��b��>�;3=�[b��6�8Y EK�&#�[�2���g�y�}'4�,.W�o�*�,U
��P�M�+"z|��f�
6�1��d��p@�c�]#�6�`|\&�腗�|��q(neH͈l�.!�V��!���G�0��W�ӓt�����
Z.�s����ǎ�J;��������p_n�T^���h�i�B|����7��;���%���F�/�M`�N�)�I�=����l�r�Y����Y�p��ӗ�ŋ��ӽ�@N���PF��S]�֧�y�CI��lico��&�n/W~�����9�9���j�h���4/��`;$f�J�I���qWH��f�ƅ� +[$�\o��f[�SK�k{K#o@zi��5~R2��!p�b}��u`%PEZ�?s=�;��_���$��ݴU��)o<.�Ng��7]�'U�|�w0�K����j�]v>��^K�+�@�@�Y�U}�C;ƗS>H��<�K �.ֿ���p�D�B zl�y�w,n:�dcf��+�'�;���]i��4Q���|��!@0E�;gwKE��Q�JHMM��<�B.*�ۛj��el�uJf���D��LsV��_�>5�r(�Uf�n>_�����?5)��e��l��Y.Ao�"5N��D�&�Ѵ G�	�&��������G�5,��>��I}���"��ma��=C���U�)�ފ�)k�N�Cf2�W₴��d.Q\~NE�� �'��o*>�؂�v�;:�Z�^Zm�V�(k���ma��yF�*2���Z��� ���(��/K��T�����n<�!��φ�%��Ii�a�AX��?���F[�����`=3��dJ6�J�W�1���6ݔ=��Z�C��>���5т�5��䖭o��?��inݲ@	E�6�G)QR?^���>:�;1~:8|LJŚ�n��C�S��\�D���K�9v�2}V�6�GQ�¨uE�#�Ø1����>V0��es|C�i0����] N[��6��8�;A�\�|S�d9��vs1�ֻ;Ve��i�Q$�@	��b����#�y� ��l�H��"��h�v\�G���>�)Z 
�G6�zП&���b������v0�����@��=�
O�E!0w�!%2�$��J��W(ooH|��%b���JBO.J�̠�I�� 2���i�@_葅�M�� 	�ac�ҧ曈����ƮV3Pg�ȇA�x34Č _W��b7��u�j��94e��f�Ȟ�<�ғ	P PT6� 9��Q7�y�C�j:��@GXd�=_���H��<hgޜLa�<�נn*>u��HS�HI��qw�X|
'���i�C�&Y1�$��l�2,�sJ���o�saƄ��4����~o��[a��q��71t��(�;�BX���[nR�JL�}a�r*_h�8M>��VBB��v��_]w��qצօm⟻�俦KA���f�����~G{�e����}� ����#	�/>�ᭈвf��!�)�S�=A��&�z����r2l���<�]���n1��[��$!O�3�ǘ-�I����Y����W��ıH�r>�6z���ʿ!$��0�$sT�+8���n��1��'l����ni���36��%+��
^����ߧ�L��D��k��f,
VR�OR`: �� �nm�gH��x��ۄ	AW(0�=��B��+s�w�<�*�M0Zu��5����2�'>�i��y�(�ޓ�#�G����U�߼w��,^%���"�̤��?� V���;P�g��Q��ۚ�35{�� A������E�����
���\�ַ6�^�H?�M�"��$�p0C��3�����쐶��(�j�+]�t�>����F2p����!�3)�n>�(/��K���*Ab�B��J�S,u:0��LV&�L@��/�+zt�)��Tm�ͅ�pcgN�ݝMh�L�/s_������Pq�t���;�ʻb/�J�:���ӟ� $��b��'��Ik�ٕ
�p:-���}��%��2DĴ)ks��M��Ar)���ƈ�FP�z�+)#�!f���MoᴪA��I�pD�ߑ���ď��P�h2��&9�y�O]Az�:���+)|�b=.�݃�5�Hݕ��( !&�jyL���d%����g���/��F1l�Cj��v�KX�mf�fe:{V[��p-"!}�1�3|������(��ttt��s�Oũ���!��r� �����=l�5%*ߞR`(w�l���t�U-Xkv�Zel�֊��O�s��/ '�D�CT���0��w?�ˁ��Ż¯�j�Uv}򮳺V�B��6e0���`8��W˘+bX��c=�U�~���#��F��^��߾c��=ϫv]s̭�J-�~l�st.�2O��b�Vl��+l{D	xЧ�hp-0k�8��O�٠$�Z�=�E�a��rI�Kg�6/-
�U���p�7WF��9��r��N������-y�Eā�,�lA�90mA˖��?v7OZ��d�'(�8*�4S*uB��Ҩ2�7���|���3��KAm ?c��C�����e���2*�I�m�We/_mu�(o~7S���~aّ.<���Q�8���E[>�]�����uT�Ø(L��_�N������c��[�_~=��s3��'�>d�_�P��6U!�!B��4�����&m�h��v7��_<�W��;�R�m{xr���P�-����9�@Dn�{��V�>w���R��ʁ�];�Ɠ��I�Y�d�M[6ݶ`k;���`�)�+��2��&Nt��Z����4��:�1��l�)�Ot���+c
��"뉞E>|@��Y/v����,
2�>z��;�����X�"ۼ�P��P9كR[���@x���̭f�ʞ��{�:̓n��ld7��$vv�o�^+)XqQ�'՜����>\m���7%�)��QoCB#� �ew����+uV�'�X����ϡ�Ra'���kC=L~=9�ڀo�1��v,Z1��%��A>)����R�U'���MӍ�wPFn��Qᦔ���ה�� 6�Y��t�f�d7�*�ڨ_��9�]:�8��q�	z��(���3��ѿN��i�%U����JzDe�k�i�e(�%+�'���Hߞ�`�S��A���0s�f������3��rǻ�\��|�'���w�eMd�=�3���q��L(ޯ�0^����̘fն�/YS��R����N�t	G��_���0��$XH��y����&��rJe���^v%�}i��ہm���h�|�g�l�R�:���\|6����g�&���1�ZM6��#������P�n#�,�W �rp����BW��R;����If����rJ��r�cʣY��$�O$��g3�R��ֻ))"B��K��6�C����&����˚amQqE~Lͪ������] ���K�ט���Ɔ�a�,�P^��9TM��`&ҝ8[�1���\�@�5����	��xU�4(��HA��$yT����e}"������l{?�f�;����Is��l�=�s͞���\��PV�I�c��7m�/�ꍪ��m3�ys���E� �����C6]T�MZu{��`	�g�C��߉ª�(���0ZN}�M����x3E4�؟��L
}J�0\c�/��'ȱ`(����?C��Gip�=	�P> ��_�Ţ�;WH�l�x[�c�eH�Ⱥ>����nl����杘��C랁,kf*<_��ƺ���?��6e��UY�Ӵ����18� ���o����c�6Z���%������`\�6R�ߩ���mW�Lgܕ�s���m0�.�L���7���)�B�Zls��e�~�P�S���e��C��Y���dCҁ����y��U�c4y��n@�|UB�հ��)�ژb����{`[n�)���[�Չ�K;vԵPלM�גO}�X�\��G�<�I�Y��@�T�#6d�!S�l��8>��r���q�����;J��)�\��Zh�k���e�ˮ	{	2=��E`���8_�+?b1����2��OLj�:�e�%k}�� &��*�`Ke]a C�#n����{+���ŵ�� ��_��C��P�D�׽X$C��I����|������o�#�c��JȬ��Zo��" �d�M�؍J�7�}��F�@ձ �ilT.w��a3�"�»��ơ�����Q�!�ߧƼ��-��P�]� 9�C!�e��DY/̉"�ѿ`��pc�����ͮ8?*3������q�O7a3�K]u�r�U��1?��껈��Ϫ���ڒ���$�9I����~�(�i\y�(�ř��� \?���-�v�d��h���z�9o��ZK2��r���5�q���R�J��j��kܻ�Nd����g�B�k�F�6�;�����1&8D�
A���c�!~'�K|�+^��/��p��8��}�I
� KA@��C�S���S*�%�/�'��+�:���w���������?a����fW�I>���\aO�B�E���1��fɊ�Ka�!��ɝ�hչ6�G�c���D�%
d� �R#I�SKփx((��Fl���㮅��q��K���5�Q� 2H�y���e�E lB��^��ӱm�j��v���#	�vJN�����ڟR+�Xs�	��-�z�gM��ɸ��|XC��6tP[��kpn'���U���M�����^����{y�8�V-�����-|[K9k#�X�D�,v�m�<r�e�LP�>�f���Q6��Ŷ��8A_1�v3~�8����z(LЖs�^�Hh�/v�����k5��r����yd�{�w
�T�38g�Xv��
����bo�P������Kg���>z�(r2�b��uؠ��,&&���й�*���y0�?H;��W�A���.T[�sۗ)�>����'j7c~!�qrm��ù�J��Tw�������h��$�Vӎ����y�:H��=�!]`��f��,8�9EL��i�T/5Ù�r�ޫ�w��m}�
!�$����7
��_bV�WǓz(	�0��E+�f����`�����b��i �ZY�|"�|��е#�'(%��7��v��]J���H�� �vёy�s/I3����ד���,5�k���TUG�x��U:r~J�ȅ����U�&�G��f�k���y7K�f�ؙ&l ��y� DC�B�Ő��N� �(f��㌣�6�I-��r3�x޼��� �Y�'�+F�؝ɑD�L;{.�>�ѡ��JZ��˘�U2�I�rF����P�ei������)^���X�W��f�#�x���:�^��*�,>�������#�n\��0Ӻ��F�P3yB<�%O}K���e�È��a	��u�d\�b��Y��#�|:��Oa�IB�}�	+b�^��yUV�+x��D?��B�ݩWYb�b��]S��e�������J�3zh���쮊���ħ�����@$Q��B�ѠG6��9���5���8 ]y
��(G�/��L��"���N9kϷ����q	ӣ^^�n�E�4p��h츤Y�u;̌�)��_�#ls���0����V���b{����Ң�Q^�4qk�V*� xXL��>g�桷�=�\P�S#��'�V[[�w�K���@%zFM��lZs�u��R�Ev���V�3J/Z�P�Q7Z�4EN}�*7����l�#��K=������� ��RL��;��D��	�'���+ÿ�j���s3�e�.Ҽ�T�h�R4(N�⌁����|�J*O �9]9v���y��n�mx�C������CnP_����,[V�J����I�����y�2Q! x��@Ӫϐ�Lr7LCW�ɘl`�P�kOҸ��	b)���X^xɱ5TY39�W�v���%<T3ec��}*��/�<�n|)�P'��>j9�nU�؛^Lɛ��1a��01��>�E6.�fLAV�I=5eʑ�����˵4�~Oq���/�8���r���p�}j�S"d����zR;i!nX@��"H�	v���jU�D�z5���ǝ�Lxo�C�AĎ'�*�������G���,rb#�M�����}�!O��(n�mAK^�T|�q���{Ģ�Y薥B��:�6Z���w����3s�ܐ2 N�����:V����D�E�tF\2̚�el��g�Ib(a`t�jV��YK�؋��c�D �
�,]w9�Q�bȡp[�Of�)zG����O�!���)
���N}�+�O�R�O$�{���C�}m?,�z���|M�k(��D(PW_e���������:ߧ?�wp�ۥ:�U3��xn���l��!U��-/B�c�}�(y��\:���q�X�?��X�8πWD�����lu<8�	v6r�6PW�߹ʻ��1��U�G:3Z�Ѕ1�f�kP�B�L˥ux@׉s�=��96�]��st����8�9ӛ�����ͮ.�`�4��Q��C%R%��/�����<��w7X�3�e�
翺���S�~�|���_��R����k��> ���R�o�lc���L;�`5��EӒ@]ӳ6�i^��o�b(4W��L��DF$����Sƨ���^;:N��Y;Z�X���@d�;�O���E?��!�@5�,G��� ����u(:v�?�<��Jn?7�:qe��5����2$
z�k% �`i�(���8FT��.X[f�p9�뢑�l�\��e�Ԅ�A��>�SF����������w�d�R
"�s72��ci���6mZ�:<�=���\�M���}�x����VH;���/m��M'�7�	��,��#���֪_'v&��X|q�#JN�͟ƹH��:� s�fǪt謐cvN�[��0�����R��)�!j��0&Z.����&�W���.�7�?��!�>��Y���q���Tgܘe%ü���? d��%��J���ި�KF,�a1��N�*n����`{�$5��ב�7B���R�����A#���6.�\J�PΖ�5�]8t3�'��¨A
�£�j���L�X��fuZ�fQ�@��Cop,%xV��nVL��B ��6 �!�֨%�V�j?���ؚE�F�r<��frq��V���pEdNk���ȳ�]���ɡfȦ���f���T��T,�������%\7�\Ky��H]��A� ���C��0�{^�ݮM�M��1����� �P����
4�"^U�?V�#j�'
`�����*������
��R��g�:�L?���I�fe�y�=��k����nj�����w
O��:�*�W��Ah��'�͹�̦�f�Q�Aj%���D�ҵ���ER��lH¼���s�����ٵx�x��i"��2$�E���Fj��M�Jj�Y��c	@�y�	�΍���ud�F7�\�nD�a 5��e�]~�2���5�D��|���ز`TuN�!�X����IwqJB�*~���<`+�lj��_�7,Q�)��}X�����+XU ["�v|���}H��T��6�	;�k�X&��I�u�E�ȼ�B���"8P�\���[�}��[�_������������T�0��ԟ	������v�F�/�525.(������E��B������xjS���;`6������[�b
9���P�N�������"�sh �Pq�l�2���1�����p����2��uYSMQ���E��e��H�!˻^�cP���N�mxp���p��F�;W�~-�Y�M\�S5\�{8o�3W�Y/0�7[��m/F�0=�}�~�K��?���A@@	;9�gJ��ʷJ�:,OcȔ�&'�C�w�K!�bu�)a��5�Zs3�&�-9��%����>�[/��Ѣ������G����d��S�w�"3��/_{H:@�m@J p��'���L �\*��J��Z �uB�%
�
q��)1!�I&F3���'LXO�|&��D�j�  xnD���\0I!��sp�����䕃ʀ��Ywr:W�
��}��S���@=����D���4��/ksP��4����m��5]CAj��?&3��V��	�2o$%!�9IC~`@{r�LZ���T�E(����6=�2��E�w�\8���N��{�/n/A���&O2�kI~�CC}=ߠ>�K�<��8����7����bTs£n�t�.�`���$��-����wۮ��Ү��\���%?�V�H��`�}�O�`!s�<��4����	&����Rr1�iB��n=�� F�Q��8�t2T|���o���"�VA�1ĭ�ؑ
}���BA�(�6�JhZ���*؊����'򗄻�ns�rۘ�k&�����X4������T&�p����2�	�����U`5R���u��+��w0!��&��ET(�˽���fedT~���-N��[�0ZO���Eo���M3������t�����|6k��aνL����u��e!>C��f���g�v�Z<~�Wɸ���Ȩ�94��!���^��3Y����,	�4��G���=Z�fs�h��BQ�D��!��b��Qmˎ����
r'���$B��3'��� R������GX~��kCJ��ivY����e~��쉰lN�ڜ�R�?�n3�e3Q�+C�<H�\WrT��>n��K���}� ��w��+�ۤ6.3������L�5'�Y�2q�ͼ�
��*�D�g|AA+�瑩e�h�l��*� R�Ip'���B�l����=
�����Wb�|u�$Ò�>��CyU/"ˍ������V�!�: �����g3�>�_���]<�������0�jR��$4��0�~�$���S�Ҋ���|�9�Q�gz%��j1Gd�^�[�;��K���2�$$D��Y&�1�<�b�±\���a�DLĜ�XQ��9jB�f.��s���L���ǫ�.H��JН%^���A�8���nA2o��s�R������By�m��Dг��РI�N=(;����?к��}��4��7��"��M��q����Z֜1�jt���.����:-2�j��*�B�t�d�Q�x�=D#OA�����\�2�>�N�=���Z��|�)��7?��	s����
���Bvʔ�<�d�P+��s{����=4�[� �{nMC�I�|2�N~(�ꬾ=�O�p���2z�@^ڠ��KZ�@3/�au�����hJ�?����B:u
��!Rbu_]���dv�<��S�q��#����&��#������ֻ���Y�H�i{��Y���@f�*�G�k\xO��;�UX�@ga��ڐ�Dk_5*OA��}ѹ�����S�ZR,�L��O!D2SPG�8Ք�ׁV�[$��Q�V���ǡ�=07U���4�_�E�_����Tfʿ�Ӯ���Q�80�P�&8+�Q\ۄ1ÝD�J�r�&z����z�5��:�\�� m	��, �mK�l0g�� d��'ڞs�!c[��4��0���@��+$�0LHI�z��y�~͙�D������R����%dP�t��9�YN������95�~�GXK��Z�}��r��1*v�4��{uz�0�ńAG��ճ���g��SgJDL�"$��ih�/(q�w�5�mV�M�*�LO ���ծ�-}�2����홢����g����w,��)��CuW�c]pb�	�gJ�Fq"hy�M�gX»�c8+�{�o��)��eO�T%�w���K����%1A��,��P���z0]2��t�2�V��%Q(��8Ɗ��{�dP�W 4Y��Nc�F�ҳ�xW4����� 3��P��DQiY�[��;x��������YgrT�!2l�9_�n�ˣ���pM�c=1)��u�h�Rݘ��	����g`�mC����@��â���س�O2D.F�E�RQ��̜����F*�]쮌]�X�_�Of�`H�Bi�e�ń*:��*H[������(t�R�]�;�q��m�mξ���`��eO-�{(�F����򑫥��c��d���z�!%��v\��?�B�ō�p�v.����'&���j6����+�鵺���:�Kd�4��O/��gf���sĀxh�gC��A���*��q�Y���Wʲ�IWZn�Z����'��:2A;�VK�@񽾬[��z�� A��&@�!�൭$��Vl�^�g �ma�mTL���È���)>}Mۺm�N񨷀6'�����ޢ��7�ۑ_�rR��LT�(�<*:v�֠�R�"k�������L?��d*�D��o��'�b���C Yl�F�d��� I՘��}���`H�:�Z5�i�T I]
�i�*�8*���G�nP�)���,0��(;*�u��S�u�;�h��|�Q
{	}A���rI�,��ʼ�0p\n�$�A�U��_'m�	��	�1������� K�䫊MI+nu�,��n��L�Ԯl�ã�x{RD��4�n��zAm���5rڔ��u�L�.ژ��|�q��,e����a��"��40��PD8�Pk��`��	�r
�!���OT)�Rܙտ�����'��.g,�&3���A�_@;�{7)"�&h���N��&P6�QkHEvRd@���IH�q}�WA�_���L�l�n�U�x���@�Z����ݾ�Es�m�G��\���9h`7� �\����l^�w���)ɽ6>�Ҋ;/������7���SvK��uQVh�V��rD1�/B�FbŇ �%C�<��`��_ϯ�y�Sm��J[���Mbd�j�k���w���Bg@)����ܪ˸��oy3I�38��Y�V眄"�^2yw���p�0��l��%ֱ֔�z���/%D�3�ɖӰ�V-c���a�h"%#t��4[���tH暜�1D��2�0Ls��r~������L�]q�/�y�^!����y뙎
<)�b���ǫ��:j��$<���z�|�?��Zi�;Lz�&�c���5b��r�H�+:�t~��7���jx�]4�H��M�x�� _Bq�G#�#i�F�:��r6Tq+W���u��mؿ�x�P�CjP�p���/�xˤ}�U���ei�~���8���Vg��%4�9K�=*:Q����t�wW��������<�����5�t� �ʰ���krF�g��YX���A�2��c:�w~�E��������䋪k	�XѺ���b�K�'���Y^���\,�sAu���գ}�w Δ��!�6u:1T��;"s�&*����
R�<TrC��(����{J�>����s��nTB�݊�qX7�����w�-&�u�A�Z��m�2>��G�p��4Z�E�4>j�'�;�E-��C��f��ד�-Ó����D��k|)� ��aą|��-�����A��ڈ�zao�6VǤ/QLqe��.�^�.�UQ���@�
:5Ĭ�W�]cTHÅm�W�������VI_d:�Q�,�[dK�
T�K��f��df*B���bxn�]�dP��6����f��n�a�E'�}��/�E�WU�EJ�~�Cs�E�SMPC���J��t�ܥzM�:2Ƃ�G|�8��?�m>a��tB��y�����b:�U�)Nˆ߽3�1�+~��̞1�&�pnlE�BՆ��$Z��L��/��<�*�z����H�����Ce��/2f\��<dq�樔Py���d�Q!���u���_h��`�8���|cT������#�9n݀���)�@��HNS������*����)�Y�	�������g�7��c6�)�_/8�l'k$%��t����{g\�����׳�NM��@��}�(Fl���!��p��E�V��%!=�A�
�YKm����	��3��[n��fB��׍RW���Ҋ��N�o��}j�G�'�R .� E
��-�ƅ[�~Q�G�|���y�Oټ'�`��G&����[�K�R8)#�%�.�U�
0TY�[���)�g���=#��:4�gꦩ3���vPR�|<�2�#69@?ެ�eЀi�.�����z>ֿp[�q�<�ό��ω�HBٛ�ܝ F�r����$�y��B=�0�i�_1�%IYՕЧ�HIxD�"��#��N:5���
G��
�4/�aoc�n/�2�{����"��s��#8t���/V4/�pn��l��Ƌ�x�󯋪���T��H}�.�_�s3�;�&����H�ɀ���B�b��v�s[L�K�8��D+���9�%������X���8��	n��\��3�������7���g[pr�$�Ǡ�_�X�F�1g�Nk�����?x.���*�?��E�E}�3n�'�;_G(���Q���AOZ�
)!�}B������x�^����	}�(�wz��J�%ѽAnE��f�-�o���9aK2w?�Ρ�KL��N(�A�Ӆ�_$�s\�}�R][�IZ��6�Ҙ�
�g��?;͔&#�S�k�Tu�G�v�m�vX�+��B9V�U��x]��R��l���*��J�8�!��d�@�k�l�[�:���@�aDd�*[��������v�2��Q4Ir0�m	WG�i�3h�3vv�L
 �Q�a�<]�0Y�P�.�l7�xw��\H��cR6�����4�C2P
��j!E�CX�nϘt����s��&n<�����GU�^�7��#38u�z/�T	�z��Y��
k<g%iX�ʃ��V:�ZU��v�>I.�(�-�xO����TA��'DH��	Z%;�͈}29�jcs�'UcN�6�ӛ�]q?�G{w���58��id��_�Iʯ�e�0�l9[s<����V?�\�2\���oN���S�%���'�������H��`��
Ǣ82#:'eqFo/ʦD�חfÌ��U�*oTi`��<�Y"H�e�c^5-���x^B����;�ݠX��\�
��y'%�Xc��&��+ �8��zf�����c|�T¼�K��8�I���*p��㇪b�3ۭI]�����Q�&�D�u����fL�荫'8D��1�<�vf+ӋQ%����?̬S�ą�9��mY^�!��j�å�ܺ���S�EU����R$� 9K�0�UH���nʥ��q�v����[H�P�%7YW�����l�D��Vx��N�`�'��t�F���:h��8�S^����A��ż��lw���֫FJ��!)�>U����Y�c� و�J��7_�k�Z����+V�՞mX,��D�cE��1�vxOZNl
��Q��	ԏb�@PQ�h�-���V<�B6m�T;�lC1�{�q+�mM�r���V��T��S�(	 &�Ǡ����4+��k��"�%Q��3C ���@�C�`9N1"�F�q<��BgR��z,4��!��#��MȺ~9���ŵM�� ��7�S�$L2�+��y�CL�W ��̞�� ksd�	(8ʟQ�rE�o仸� ���Aq��ի�VU=����q��륹8�r��ν���R)����n{�g��Xդ"��s�DUo�R���KG��.�{�Ԫd��f��$ė�5�����>����N���Ha�/�<��¼҆IV�D)Jr�u'K܃8��@�6��u�cC��y�>+a'�/����������7㴔��[�Ѳ���G�l���0?�1���N��i����ȝ�{?�a<��uYT�i ��g�2*��ݳ����G�Qf"����h/���||>?�c�Ab�fN+�
���	�Q*�b33�M%2���N0��'���<�k��e��pͤF�R^zK
���=�P���ك�j�lb^�d�/B��+k���G��H!�]���\%׌n���ڙ�e�?3�ˢ*��U�@��:��7,9I?��#�|y�.ה�vl=�إ|~!���D�7s��N�v��b&�5����b�L��@TG8��o�߭�wB���_�oܾ�;�I8�s��3d���jZ�#���淆�\��u>7�A��A�g^"�r@�E(�L�n����h�ޙI�X�Z]&Q�"`/c��0��OfHU��]���P�cO*�(l<�.d�L�`U�qk�qm)� �% ��\#O���3ow��Ќ\����|zN:���mV��0��`�V��L�8A��{x���lJR�n�u��K�ioX�(�4 q�;xI01�-T�����~�)sO�R�!>�-W_��-mk����Fn��yc��qKdΉMX2�`���H֏<�ڿ�����[�<������>�#;!i3(aD�w�P�"�bz�-YO�p�=7P�͓��K19�?$�CW���������$``�=���;�ZM�[F,�7���5`�\��F��`�Ng���o�}(f;2�6\!�G�G�B�O`�k��A������t2�6ݑ)�V��z�2��F혽���D�W��R|8YXX<ąp��x��S{������nM�TXeKw�����E���\w=�.�
���+sm�Xn��e(��<�%G��D�I�[��U��v�y鑚5G���� -�`-�2 |/��NK�s�Y�����M^$��Nq���+��=�)R�]���(�$P��lڨ$��.տ2����,���:\�����-�S|�%��jPPO2f���'�q'a0�-x�;^6	���Bsv,�4|Z/�l\Og*��L�ܮ?MjNR&WF�h��vWA���v6�p����\���C7ԁR�*6"4>�)%�1=y�O,�j!�4�)��:��wg�'��C�QI�廉k����k�3�=�����M3�l���X?g�n=%�k�q> ����I����D�8,�7�!������������!.�~���$��)v�u�{7��/'q_���x ���q�GU�ǥ���l|Գ�M����1F�ăW�-k�u#���o�O��W�%� 競��)!ē=ԕ k�H�1���נ�8����h�k��{o�!���B��g6�`��o����H/	�{�ھ;H�q�� [C���s'@@�kf��������}eд,��H�`��;�c�}^�I\���f�?�[h�L���Q�$��VH�P����/��>Zs����t��Cp	����b�cbpz��`��4�l,��76�y��Y�@�ɴ��ڥ ���o�����DN�K�Dlw����:�(�g���q���;�#ָ�d���[�G�3�Al��ⴘ�`M��L<J�@ǘ�����F��� ¾y��x٫�E%�Yݮ0 ]��ܻ�1�&��Ѫ>��}"(;ɔg��vق����tiq4d�)w���+XF�h�'	���o/I�s�9����L=�8"gA׫i���$&A�߈[��� ���w�[3�U�M�Xij�q3�d0�9���]e~�J�b�&!=G�a�|lw�-�`U=�����t5�G�bq���ê�CI�p���+/,1�}CUd1m]S
 7�(��2������؏�Zd�r~�ҫ�;b���/�x(���`���7kUg��HcR�劌��wP�5��}�L@S�rp9��؜��ah/��E�2�ü;�3���3�K���UMz���!���%��O��2��a��v{�����h�]Nw��*Ĳ#�낺����p[>l8���q�?z�����u�\o7]�jF�L�?�w�5���w���2����#�Sn�Ue��z���}A�"r>���|eP���!�����2힆�r�á9�*Gv��Hڏ�^�]��dvIh��J��Q4��&{��l)G������q���v��#�+��cv��n:Į��?b��t���PBۇ�	��;@�P���/o>1MK�c����3����K�(ЩN%���8p�t��rr���WJ�X�J�QO��ԅ����D�;�Z�l������Rj�,�׼�΢���=?�+���l�;���xm:,�������� h*��w
��Yh|���
�6vu��;'�ް�n=/�����)�w���'H,���6��	�Ci��d� �_�Q0V���&5� Tj�{��h�"I�E�sq,8����=[���yD��S���Rg�LG�ǋ?��}� �Y5l'@rQ4X�q����o �A�g9{���K���jF;�1����|ӪK�x�Iƶ�CFxsv �b��a˩w�f�|
�V�1"0�2��k��4m��'��׈>���׾����)�G�In@hM*ۏށ��V/AZ�G8���U���ʤX����7A/xኟ-8.�c7�g��/T*T2�?��u��`|}�+�K@��O� P�	g �������z1fm�+4�YZȒ��z(g��Z�����Еyž1�ڊ5��"C�M|щN�K�&���=�0��7C5������W���W��e��-| S]�阮XYf�R����Tb��E{�t��Nb�h�U�ŧ1�Ͼ��Oc)�&���L�"J���m絭"�ڼ��_�+��Zhu .�D�=(����Xe�`��ޣO��n����L�mb�H����6v�c	P1��'�x� ��w����y_N��{���]pw���3,����<�[\)�JS�8q��#�z���	C�Zl�r1�� ��8C�v�x}��{ܺ0^�5e����c���[�A�	t����$�&�Là5-h�M����X�>��`���Q����ɍ�~��VOz��/�DA݅��O�(��P�2�$_�#.Z�$%���t �O�G�8b�T���P���T��"�]�R�m��e� ��K0R{�f������1�#�7LL�U�+h����h@�9<��ZYZ�G!���Lhh���=P$�9X��ԝ�H��5���Z�t�G�Z�8y���Rօ�c���B�/��U��ɤ���sYT����s�anX�1kQ���*��<��W.�� +6i��v4�5:"dyx��O&˨*��8�s^�]U���'�Mgg��]6����4M�\q�Ƽ�Zb�+ �:������,']`f0�;��0��d�W������Ky����uԘ!�e����)�t�ಡ��~�$[��(*	Du� l"��0m�6���T��� ɟ���'��?!g����J� ���*s�;�v|$�Rh/���"��k�j��<e�����/v*���Ĭ��7�c�,���Zi����ڙ=��;�����g���ѥ���\�>��a>2C*�ĽW����7��N8�2�i��׾�~�_e7���'$���d�s~��جOP�T�5�ڳ�+��mY�����Lcu�����P�1�IWZG?l)��M��t� ��90h��^���f	"�����4]��
�5m��c��IVz��
��c� �_����p�X� �Y��O�M~������/���zZ9��c¦ȖB��ϹZTD<���I�8U:���{��o�O���v���ٱ�����L�_[
P+��n��?����w�� ։S�t hG� �Uߘ��dڶ �]�V��2���u8�h?{�PMM�A�\�M7m!�0�i���?��<&П �+8o�>�I�2n��P���E6��$���-ig����n�7��g&|���h)��+-���L�A�����-��	@���P���7
J��Go�ڳ9L��f-�S������#��˴�ss2���|T�#��De���bzK(Bܔ\Fv��^�8.��E��NB�Ϝ�j϶>x��xl�|]���-L�=冸���ؿq��-�*۟����������@ \4b�x����|���:��R�/�D�Ks��\`��|xX���_p����m�,���N�m�	�u�'؝=����'�������} ,P����^�����aG���e���Yo���G9��Ryq��D��4�}���[�bn!�����Lq>לy��:f�����v��uR7�R"�>�|��>���0~��7����X��4�A���\���gݹ���x���37iD}�"Z��Խ���ݩ�(5���DYPѦŷ���a���E�SB��5Űf����@f[��7�(P�	f�౱b\��{I�	'H^�iĠ ���PB��%����1�"lM19�4e6S���g�i�]��I�:GV�Ė�z���vl�k(L}-��auD,)[�/�����#V���RE7ϸ`�J_R�f�/sM���^��χR2%gyǗ�0�7?'��~5}N����h:�V�c��7��z��o|�ő�Lp��C��4LIm�q
_�2,�]�`�8��8�]7��3Ww�a�X	��Q�٭�64
������q"�n�!�tJ����.�H_�*�8�@�׼��[I�(~�s5��c�	~��/���4$L�B����ˉ����O%�zB}��CV��W��L�����zD��)���������N��g�q\�Z���6���2*�� 	s~:���@'
�!���i��B��e�d�T��:�Г�l�<AY��jX���{��'-�q� .c�Z�!Y����<q��4��rm�|�R�UO��}@}�o�HS��h��@r^�m���%BXY��plݲH�c⾂s^��8̊��~E�dZWgK��f��m�i99�L�P
ZǤh׵��
8�!�� ��}��"CpzվV�s	�o��NqO\K�B�Y�P�9�H������?����7?�X�*UJKWH0b�/�a�����W
g���=���pC\�uC�;:g���Y�.&/vO�@���W��&qY���b�A���n����@�G}�yx=������$��'
�o�-��QΒC�&�t|���e���+_!���ê6s�2���{cଦ.��Z�+I�k?�U�I�����]������y�lJŸs$꣪��}A��X�?�]����p�Ћ��.깕���u�AՊ��W���4���d��h��������;L�ˇBڤ�v���L�DRb(�Ju�A'+�<����4����*�±���]�m����Aa' #���^�`~�j���j/M��&�'��a<y�kB�$鯵h��D<?�˟"�{	ˣM�y��7K�K��2&H��9%|�'6��(�"	�<BU�K����ș�,**�:�+*:	Ɗ��جr����i���Ց�;p�c��d��@�eΜ�����3��F��	�g�
����i;+���c�@_T��nu�x�T�<7C�v���wZ�W9tF�4��4���O�9���,e�ѼSx�g'�D�h�M9xW	��6��I	c�u��R�>�&�����,\�$��ZL�D*���� IX�=�%<���t�9N������nor�WM��73�8`]l�~_����1,�!z�ѫ��u��Q�g{JElJ�U�z���E�kÍn:�aN�X>�'�*pW�,��+i��PYڌ@������j�T�C�]S���z�4��3��d�%�x$5�UӍ��eT��	Y��9F��
����B1Th���\�6р�l7��(������V���m���˪|�SvJDir�/I�gj@$�=dKY��c����d�����R�0�=>+�nZ���G��B�I!��7���$h���S���R@^�4#�f�D���<��mU`�Ê�JΜ�2~�0���������ZUd��?3��ѧX.6K����[��L�m�&p��d\ to�r�o!�+!��(����|��E�L^۪�q.�'Wk,��]��U>���(�u}]WPO��U!���aP����^�G�8!��f���jB$9v H��y�C��3�k��Y�?E�P�ws�.#�=F!�->S(����.b��I��H��g���뜕�=T<��Ư���*��j��\�����Ux�Y^X�{����9ie|ǁ�g����u�OJP�T�m�>܃^�.�ZE�b��� �$b��&ZUT,�y���������v�A=	��������N��-�LvzS�R�.���Y#v�H�#�}�� ��_b���^�r�&f�-i����,���ҥR�ԁIE�)��wJ(?�5����D��QXc���]��_�h��+�����MM��,��[2��Í�,���s�3���� m��Sĺ�@M��
�I��ɹY�EO���y#�z �R�� ����D.�W�GΪ��cc���a�9����%k������yzp��IH�$�xQ��(�g��{V:B����_�|����*�ߠ/���|� 3��Ы�!�M��)2���fDB0��Y�}����Ӊs���b0�(]"�t�xU�����<�����l1L�7����'[� ��R�%�H�����S���r��u�.0-��2ۧ���̶I�f���u�����D�'9�����������I}��{�3�N�D	�uu��q�	 an+�}��@�$�(��G��෨���>)J��#��*|��m���xD��D�1Q����V���(k���Qi@k֜����@ r���b�2"I`5��@'Õ��{L��]�<��[cfH�U�̺?�<�"+�2�1����P5q�!@��� �!�n���q��wpRVx�@���Q!>j6���7YF�7�?��Q�����:
�_+�3��
d

`o�ۯ���*<��=n�m�戇��%�	9�"�Is�V��e��ɝ���wr��rĿrU���Mxڎ5�6HX���=��S�>1����~�VH�f+��X�l�p�Q:��!q�&��U�^�*�cv�xi���4��YfAaWG��/�5�����ms���Q3�����W��'���vFK����yU���ϻ���N>�:�B,�x~z��������$�!��m+E�Y�-���v��6j�}t�h�Y�<��9������$v%2]~�ZV=0ܘ��c[���r�W\<����1�چ�e�ש����Vv4%H�ir�;��0�k��� /s����^ػ�YQ���1TI�Ќ�x��J!�=�4~�	W���n��͈U�p�.����c~�2���D����(�˃c���\e�h�R��hY��h]��S���	�H�Q/xrڐ��Bq�=����J�QU�����?��Kg�ekڔ���]7}���� rTg�X��H@g�W������Ջ��
Oe���SA���_]����>�|},�i�X#�H�\=۸ҵf�3q�0?����+�K�m�
!�<��`���{��ܛn������閾;M��7����$oI�i��&O)?�!߲��m��(����&Ѐ)VZ�$��8��P�2W+4��ǡ7(jA;�(�ksE"��fJ��ej�O2��R�kn�h5����^�Qd-�}�	FO)-�:�۬�)��V�����À:മe��h��@$���v�?���4�7<5lW�� µэ�EfK2����:���!h2	����ld�f7�_O��]��f?~��_�֕a8�g.KS$����p�<��=f�CKCE���wBQLx���s��\t6Ҁ�h54|WR�a��u9���F���_IT]�S>Z��͐Sv��W��������FdX�6�@r����σ��m!yq�P�S��_%	�5�Rx�h*���y�U�$�Kc#�C���	����_���r��#'v��KG�\W���t��*5���p�/&�rt�x�Bp�ax�!u�+$;4C���I��%��'p����y}!G�⍃���gR!M%��ZP�T.sҀ�[���q@�]����-Ƌ< ]h��Sʟ���Vt����N;�_J�����;�M�EԲNn��0���%r�%�C�.c_�m�L"��� �~Ka�N�
�Φ���w�q��֜"���Y�\�u��r�@L_�	�'�n��xﴤr3���'2�
���%�3����rDu�����k"��Ub�{�K�d��u1+T�N�8�??"���~���+[�We�2���j�_1'�|�~��	U^���Ј\kPy7�줶��ʴ�"��OGw�F΅����5��rcBu�x���d܋�=��I�.m����Bkv&��?"�q"ؑ���m�%3:�Ѷ� zU3�J�����]�U�M3BHn�JB_V�z3���K9��c
T3�a�C�ȨƷ'���e,����e^�k�V�gsM�g����[[
�����f�5�<i�U��T/�"�ky`+����d��X�F� �cUb���s;����,&(|���6������Q��?�^�_�0v�׫�:�ZD�PK�;�_&Z��S�G��'�d߬��ez	��/�C��� s|+q�d�Sw�T��b5�ç���1D�v,v�)��S�:*;}i�h_�h�ܔI=ޠ� e��v�|�+ �&k6��dƦ�g���b�.� ��A[C�V)�b�|MG���|T>?������rp4�XQy�����ՙ*^�8�)����N�M�1��X�����Ϟ�ḫ�*\4��ʟ{�PQ8�z,j��f�V�}f�͎p�S�M�%q��d��'��N�/�|���œ��r/Lܵ���hS���tJ�]i�:��k3��7������(�/�0z�i¸�y�>����oh���jK�5��R����"�x�Fc*F���Ek9��댹+Ϥ��+"5�/�������O�(�դPKD�1?��	 �P�e����(= .��Hi[���Q�����ܷ#�$xvT�����ܯ�&���ͭN��1�,�~��Nf�;�V "J�:�Frb ��:TB�1�����Fq�x�nd��K�y��Y3��9F���Q�[�Ұ�����G�{܇�8t��(_��3��!�����e��>�k���ĕ�k��km�3����|$�������
J�C]c]f1r��B2���C�~���:y���p��[�y@�ܴ?��,F��>�D�Ҭ��Q��3�3�xd���滔|b^{�����>� ��W��>Ny����fz������d��O�г��K����
��s&e�8g	ՁR�g�߳�	 �l��4K����S��x�<���(�\�X��&!C?:cϦ}1�o���/v�GCd2K��ةU�
�qK 5"{7
�E����V�E���&l^���4�3�3�O�n(Ā�)�t"��R�p���0�YXJ��r~xie����B���2,<ȶW���5��b��*�
%�J06|��[S�=ul��:@	K\�s�U�ug��ZU����{�x2D�{��+�p�N�h�-�N^�$RUI3>����IeR��a�'W�a���U���M�q��Κw%\3�"��3ʘt0|���1k6�b��k�v�v����y#�%n=O�}!�^vU�;��jRd`vZ��.U�Т�rv�d���+)���HM�m=1�%V��C�(�����:}��%����x$�:��5aֈY]d4���A֊��<�9<Fm��m�dA'Ǚ�w4�e�k��R�Be�gl�bͬ��{'79���9��&c�?66f{��&��"��lw�2��_r�F��������s�,h#^�S�������~���o�&[V�bx۵�U<I�4�8x*�� j}0�D=5G&�]9x.}�`��ţ�I��;�:Xd^l�Ǳ�T`��"�L�F�߻�SK}�W���d��+���&��UӚ��g�����Y�3�b���,�c���@ލC��?���`�9�y8��cGzS�i����t���q����.��ϥ��ɻ��2	ǽ���jSm�z �@z��;5iV�3tj�b���`w��iڊ/��%t�d�x5�{V2��#�_�����~�(�o޼�T'�.H%�gL�����k�&/إ����±~��+���ȩa�(�K�;~<�����(�fi�`g&�xsY�|���A�0����h� ߈U�^�+e�R���y�M+$�`��*s��f�>�.l�NI-��K6p����^�YN�_ytq�x���v���e�?�rwXv��P��ҳ��5���í0�5y�Q������:���T�_u^�3��,d��� �5x擙�p6�ƺ�\O�Q��jڻ)_�:DЦl.�*kjgΥF<�l�Rf`w�+��6��m{_��2WJ#��ԅ�h ���!{oC$*oȆނ�����O�eqmN��F�F��J�fY��pL�Ԋ�8Hk6�'��Q�*E��Z�h^��_��*���V �Ur6�e�) �7���:l����d������m8=R�Cf�T�T]X�l�=����9�~V���/������fD?�c�� Mы�[5埦�V�P

eD}u`Ѣ�e����Ch��؊I��M^���s�	1yt*�b��5��kA8�
�3��";S��2��,����y���I0��&QUj�b�mW�9�MJ���j�2�h_ɳ �7ڞ~��n��%M��MG
pX���p\m�:
�(��}+p���Np���Z ��$!�]�A��w����Z�	>K>'~�O��8�"e<�8I�i
AQz�����$c���Ua�-T�v�t��S8װ�n!rߊ��=E�LBr	��ƹ��N�%�`�臔2
�]�ю��$��S�W�5_�n���4���|Dկ�S{M���(j����I��D4 �/�`
O��֨��#m�*�?��(fq��Ѧ�y	0��7V���©��xDH)0R�8���j���¨�օ�>QYS���Փ���,�o��Xq��Ժ{**����:�d[M�Z\���!�s��:Z2�݀�D�<1��,v���*F��
��%��A��
�/������#�$�D �M�j| ��=������$�����l�,*3Ftԧ!s�:���9��#a?��J���;����,�A��(1��4��� t��U��oY�*�fz��h2\ڌ>@W�o8p�?cm��C1�Cfx�B����D�?�x�YC��D1��z��?j�XH?�LĩS��b�v8����d��ć�}�C��.�2��e�D�e�Vc����nI���Zzs5�o�B^�@�ðV�y�q1�[�VdWp�����ē�o��9D�q�v���%׼�:�++@"h�+��k��5��ɭ&�J���s5��z�I�N��IW�
�p��3�3��z�'{p���'Z*�#��R���Xom"j���C8�㲐礅_.V�d��^zZ�!%x�����)Gch�JVs�ܥ0&�&}�jX���Cbfzݢ����Up�{i�.��ɠ��(w�V�w�����Ι�B������8�ڃ��W�r��̏�Y��e�*ݡ��'CW�g�:�>�,���x��$�}�"+��S+v�m�hwkX����wX_�����Ӷ:FfA��x`\"X����v-q�ɲ�(�R��	
"�tT���W�lh�ƈOQ��p�)�"�=������lA�����9�����9�T~	т0͋Ab��K#�E}��%z���Q��|��c�BZ�;.��]���͝��{��/���^О׈D��d�,�1*�έs�'��}t)�K�_+�Cql;��f�j$�1�W�G�L��^P�}�.�� s��4�R���#�|���P7�[ʒ|�����D�D�R)沪j�_��V����PM���Fp/� v�85����ur��l�pP����k�S4Uy=���]ED���h��!��Q�P�$���ݒx�3�k��2p>d��4��YGY�up'�oMG���PR��f���������U��5�Ij��h�X�>-n�2�.��Z��/�ٲ7�d�q��R�æķ�h1��P��nc=K*�ѫ�Ge[i���iO�-
��\B_X����f�_����됸�jם����<q��XL� go*b�7��'K�2�	��dD"6p��i�.;տ��(ϺP<s��=/�)����j0{U[~��F��ᆃ�4�V���r࣍W����a�8N�]k��<�i�:���q����g*F>OQl�̯�2[���:r��Y��Zu�>2˅�c\]=�Ӻ���N���Z}��@#����2��5E����Bba^���or�i��	��0GHR{'����wFUeA��,���'scTE
ʵ$�����E^R@�L�_����4����p�_oeY���K��º���̔�lQ�+>���Ŷ����&8�n�<�|�}��s��$a#kM���BLY(�k���g��r�U�������=�� 3UU��}���;.��.g�F��AT�#� �a}
��?<2�����-��T(�l�q����� �4�0���Tȸ>H�#.כӋ��η^�h�Ց՘������r�>��iՕ��l�hw�ܓ,W�����K�~�<�u�Qx�������w&
���0�z�QX]����oI� ;�͐�TRy`����{v-�}�u"o�Sڝᮗ�@��x/[�bj���3j,l�e���=����A�Wsp�Tj�;�D
/�?/Q8{����=�d��(h��@��v:B ���#�{�)�5�|�v7���K�l'��f�da��o���0(�[M�hUbK�z͟��]�oVjN�x�d=mu�ZE$��u�)�k�O�p���ݝ�QsW��)�9R��1��S�3l�d�%��$N�������F��a�R�8{Ԥs�z= �$�v��N�����!S�J?�b�P��*̙�-i��Фt�A�ͮa�|Ǆ���{�D1.�t������Rf
23V�����1O2	~ᛈu��t���E:��K��U��AY�!�/�u�/V����U��'|��w�y�|����5nc�"����z�M���Qͳ�Yv���ZN0�I�"t8�W7�v�zB͙�fA�bb�֊���׼����
n8���Q��[� 
���E����0RN;|3�&��󹻝1���,��b�'ϴ��o�j�=�3�f�S>繇���-�#CP�ʂ����FN�a۬q�����ŁJ���GX��5s�g¯}x����v��׃��j:��;��BO�?LW�����9
�,(	�� M�9�u;�����-Ǯe	DwW�c��EZ���J��8���A�� ��^�� i�fk������h`w}8�k¶�Y�d1�#���ށ�"��`^�˟a�@QS�m���o��:��L�if�f��^�-R��׏�ϰ��w�ЋM�h~�M6}�V���}��W������SM9g/���)�Y�2h���t�+���3�T� m�����j�z2��]��1��`��{GK���
�
ՓU�i��(�DQh��I#m+���M�'���Fr���L��P!�X�>��R?��@���ɲ|r���Ϫj��xX�������S"�ǇS]�FZ���{-ҥB�i���m�){�Vf��|q�R"!s*~�NɈ����B��土�B+����^b�L7��V�+��j�X��t�zi����?g��2:��A��ʉ�=��`6���T%��5_���vk�{1R)���z�%��ޢ�H���U"��.^K���5��y�����A�0]�ӂ{� ���D���5]���I���c��'����,
՟�c<���/�ؠ���x�fI�P�����؁�0'B��ڞB�ewI�۫�SȺ۸��t�;��Ά��HxC�04PyI�����0 j�+3i��joM _+�@�E���;-�@��[O��թ��,�Z�#�� �7i�P5����� ۫"��h�8Rs�YQ�	�wH����nJKt��p���~���������q�%E�����T��^�٭�J��)'���'A|�] Q�\Jٯ|���m)׏2�}/=ۿ)��Z1���m��3&<fSyV�Z��B�`d����J�P��5��3�L_������>.;������&�:��%���"�kt1IY�^b�]N����~H$���b��~��rkv;!��s����?J���k�M3�Ӆ�Z�����-g�D�����Z^x�
7�d�M�3D� {�ީT�7B�V��gV�>.V��H�M�"\5@?���YqvE����t����*ذ͚g�F�F�6]�8��@ʇ1�Z������N�*���<P�,�8������1���`��k|�=nd'|����.�z���k&lp�T?䤷���7謕�h�����l#ҿgt��P|\Y��Uo<�{�K��#(`��/� �-]�ŵ��2u�ڔ�'%J������Y�Yѧ8S�
�v���K��������k��ې
�P)��y;mŚ<�B����H�Z���Z8�aJxc���J~���q���FQ�j% s(�4bU�������E�
!�ʎ(¯�?r��x%}3p7{�u��l���8@�Bzւ�_澌&CU�C2�E��2{�C�K��eg�XG�`k�\�W�U�Ch�\�˟�s��1�����ƿr�IU����R`�cdE�Nx=����{<$`ˑ����dh����2�����A�©�4��0*���_��K.o��CX|��;C�L�6�M ��~�k0x���R�������$?����;�A�w�cjtl�d���H��8V	������Ym�S�W���=2�!{#M��h��W `2���:��t� s�<.��qR)�Ԁ�e\�+&Q$�)Fv���ˮS�r~�3|�<�(�@s/���^�ժI���u�x�qiK͚�b�'ǎ,;���439F%�f8,���_����1��dII���[�[�hU���C��һ��S^n��~wR��
*OŽU��{)�Z�������t!��!Z>����6ZBJͱ��	Yc"Cΰ�	5�ڨ�ˠP!`fp^;X�Zg��c2�A@���A4�3�c
}���okM�+��j`�d ��ؖ���b�����7�!N=A�;"�MW��-7�x�}נ�ʂiW�yr���0�D� q٭Dk���.K������= &����&|�O������'=8���3�Õ-i�
�Ƞj�̱�[�^4��Ah��\�X��B��^%�ͩ���qQ��c�Vr*�A�XܗX_�����,T��i��/ �7�{�����W3o3�e���$z�Z��6���a�hg�S.�9�G��V�Tύ.�����O�i�Rv*�}u� U-
�mP$��BƟ�=�K��!V�R�s}K�'|��#eZ��o�%��Q$���D�˲fH�s?F8`A��D%[&��c�'�W��s�0X�Ԡ���O2���.hOe��r[L�^�!~}ǛRi��B4�<���ni�$�B��z��u�me%(�^@�L�j�����D�=�.�XX��]ϡ4�&4��n�ͱȨ�v9j��Q567#�fQ�y}NOR����w
���O���o��8vc���]�D��ל-�i�5��;��D�ߒ[[�7 b}��}��
��<Y+,]@ͦ�B_k��!N��a�Έ�8�Z(�h��#�j東���j.V����D|Y;P�P�]��X����%ِ�i.���pN�I��2��.-ʢ@#��~�r��lF�z]7�2<�3L<6�#֡ y��'�1H��Ӛ�/��?w��,~I}w����ɳ{��.�k%�'>�$�
�xY �>�g��I!ޱ�h����������+��Ƃ�q����uJ�S2yL$L���+�DK>EA��@�30srۧ���6l-L����k�7��#S��DPN�ɩ���$(R74��H����a�,�ǫ�ⳋޯ��I���ϓU�
��w�h�Q��}E����?8�E�ͤU-�؊�0�����X���Ƈ������_�l����7���F �"l�П;7�bR>�i���r�ꢙ��a�2�M���٫��3�
�C�8Ƒ`�z��o]$U�]�}�3?��n�Ӟ"��-��)p�p��~���M�nH5*o�Rr�O��wa��%Y(�#%ǵ��#*r�����ȠCS���J�O�����ʠv�2�Z��u��O�t)���A_�EE�=�F�� 
�N�6�-4��>���ߝM�n���"ְ1v��x��IE�$�.+MJDn�V�����8���ђ�"M����.RD٬Ԡx������А~��"�~��p�BrgIE�jŴ@��V����Ch���i���R%q��<V*i5�´�y~���gՑ�k�]cyV��t"�W����)W(��1��Ǵ4kT�^����ś�� g���j��byS�H�=UY��{qo��z���-�>Ci6��1c��֐�"��\�EPkG�y���H��������.t�m�Г�|HB<�KIR��`0�'?7�nƋ�'Ж�".�20ҽI{.��!Pp�
>º�K���(qO�'?Ӧ�R>_���p�s�EZ���گ	�A�����jD��^���+c-����5�iq=��n�#�n�f�9r�_3{�o]#:�#��@��"h�K����O�lMɨ�;�EA��˳�]��Pn��\]̂xf�L
~�4ߍ�Z!�\O�m�y�v���Hl�7?�EM�¹X=h���|���&��&�_���3v�"�55F�ұ��S�-w:�ِ�B$L`ۡ����yۣ�}NSX�X8�Y�*-:���|bQY8NZ�Z��PLM���6��K*���GN�ֽ j_��z�b0��w�R�7�ikQy��qRb�\M��N��e{��* �J#�E/�$��������H��3�r���w�P�G��⛞�KM��!�J�B��6*M�G��o���Fr6�Vm4�u��~J�ο����iO��WJ��o��/�9#��r4?��NA����z!<�[�KP���h��MjҤ��.��x��Ω�/0%��mڠ������zk���M_���o��n��Q�E���u©}f��TP}�48�[�<#��J�������B}hIaD_�q�E�	F�B�f�E���v���qAK	�6O��;�+CE�H_�a�e˃i�HI�f I�m��3\��`��Kn�g*�g���p���G
�c�I��J�7eΎ!;50�\�EI>��������ʹ㖳�@��iU�v$��4����(��Y�3p.��$�eZ�E|�{w% �2mM���U�[	�2X\O�vz��d���1-��Sa�ҥ�]���c̈P��fIH���U;�/Qa��`��ѽL��X��_E��޴�u[tn�ǟ�&��$�åtr���X!v`��W��3)�HP�z<8��z^�׺c����˹�z�K����9c�T!�Џt�K��5�I�o�@�޻�3$���ȣ\e���ڎ���+u���\��%�ԇ�
e�b�z-%B����5�Y�!wLe��HXq�3�:լ��O`"
�^�����UIZ���ΏY�C!;yf��$o����3+NcBs���'��/U�@���SP�D���I����l��]�Ø+�~��N?�^��3�AB�	}���2։�˼��}}j�1s�+���7�U@Ż�5�栽��������_�k��OT�Ф�
G�cy �2PbJ/���c�>Fz-��R�!��^�Z���z��`�;�ç�USP�VӢ�n�M���A��e��"~,�d�<)��*{:\&˳/̖��J��I��"`*�b2k�}p�V�0�+	���C�wM����h��*�Z���SI�J��sR��'tp{���:?�BB��~C�nZ���}��A7���.`�PQ�0�#"!2���Ѹ0�*��g��s���hHP1��G�Gi�V��ls��H����dF��N�Fy|]}�%�0U�`%�ӎZ�eu&*c*f�(y���6V9��+cJ<1Y�o���X�CUE`�B���>5�?�تI�����D�s�h8��41#y ���hi�x
�R���x���8��S�( ^ �?��O\ģ�*<��ԡZ%�B-���na�G��t����k�J>u�5�.sEuӣ?��׀�x��V�{�P��i��T����yj
p��&��c���/��?�G3�-}�@@��Dm~0ɭ?��Kxf��	�|m>,wCE	/�8�8�7�WoV�-R�a�	bG��Gz+ �H�!�����������x�w��ռ��Z=.��Dt�䠸�~�7��8��D����3=^�O)�>�+�H_�ck�ƛ�/>~`g}ӄ+���q�`��X����j��[�� �E?���ޓ��m��K�ZQ9���.5,�vƣ�D9�7>¢^�%}�Q�`	G��!��vK�4a�0�*V#)S���'�$��'���,�W��UQ�����E������j�:����?d���
�-+�Tq��U�jm�u�X1^�N�C�w �>�|T��c?Y)j���Ȗ�������֊0�SB*�7�~9�%��k��������H}����7�I��t2�*Ŕ}`r'�9�^�����"��d�:fΌe���(R:'�����/�8��D�S,��A�������Z�0���U�Eə)���'�2�k&�0[8T�gIm5�v>m_��2�8�4;�3}
��F�ꏴ�tp�K;8����[�w;�T�2Td,��x���g���/�2�*f ��4n�-��tWO���&�j:�,����>�j�33#T$+e-$���<�a0O�����g:�M�]�2�!����dO���@�QwgCx?����F3I[�����v��=Kb��2I6Q6��䅫��%,2EP�Ry�ۯR���he�C���7t��v歩��*S�R����o`V��B�5�5.�Fz�m}����KN1��T�(q�j��;V���-�IXӔ
�E^B�MN`�-JU?��������K���I�[`�:}w#����T�E t���Vi�Đ#&�3�� "h'�ѽ����[��(S(���Sy������ԗ�kԹ`XbCK�)�Fk�0�h �w/�� �H%���D�Np�[�N�'��nEn���jI�U,���Y�j�����H{b[��t#>Xc2��c�<]-Xuncph5��Sd�[s����:�q�y�'�-�w�0��y�Lq�� ��+:��Ԏ�P�hz_�~��4<�cbK�y��F	��'@���!G6"G�g'd��6�Db�sl�x��iȹ|3�|�&��N�:?�Ȣ�
��W�E�}[7-q���i�&�F���)�).����OH����ȣ׻���q0P�K��+�����N���2� [�&+zE^R��P˗�^�A�0K,VT�N)�[nO��R ٵ`�_K��4����nl .5�B�ڮK1*M�u�����x���P`[V�}A����"�$�ϊZo�+�3v�8BP�����+{��t rϙp����Q�pR�9~��w~�a�&N1y�ƻ=���\;Q
S+��6���������C�V �=�n/@���i�R�h�7T�ŷZ]@���쎘�yr4��q`5���{�FK*���ya��ه���=�'���ث�x�~Ө��Z�e�����bC��X�o���Q�jFx�Z�����vR�X����wE*ȏF�����8�%��(���Ts�W�OԳ:�Ta^hs,Up ����V��(����'4��(�_������?� �gD1<RQ�X�L��G���)��u���nR��E����k�AD��2�j�2���Y�1im�$2�V_�׹��\3F&mAp/r����\�6�o ! [�W��D�������/��#�/g�����1��4�U�^����i6��G�Ն�65:��;i����A��n�\��@����	{«�#�.v�R=L�1$r�v2L�A=W�)RBU0�3_^�XD#v��-hNX]"�'�>�2�e�J-���Fy����d�u���b���nZ}��'�{[�f����(Gɾ��NT7����FA*����*�8U��}l�9.({p2�ΨO��>֨�*�@H�)�5HĔ".�Aׅ�z�����uW�FQ�VlQe���K©:�L���{���wⓃ��Y�l�i6U)������_��E����~�������괄?���q_R�'�CuJ�hsF�'-�B�Z.XΖm�#�g'x{��������Nz��-6�/��c_U�E�R@����)|3�dۮ'mu�^�3&�W����B��EH1�w��YD�rP,����8�T�	J ���XrP#�mCI��zS�{i�vX��j�6kvKu��O�7啵����1��rb���6��i�G_�&t�(+���hL���$��ronDqp"%�	MC�\z�^�x;��[{层g�,�8Z N�"U�an�:<S�C���qoW<�əd��*�È �h�!�1�ȴ����0x���f���96xun�}�0p�|�'u���j,+nc��DU�^ʣ��<�w�_L`M��n�a��L�)	���:�����̤ R��R�&�C�=��y�d��^����y�yW��%� ��2.��n�B�֪Y-�մ:�_퀾1��[�"z��y��b��ZT �Fn:��M}�t��
������/���We=��ƅ��d<U�dDX�[�jl�܈;�-���<LW߉�Z�R^���r���j��Jn�Bߞ����<<�o�<4us��n`c�Vp� d���x� �Y���L�ϼ���v�%h�-�1����,	@l��x+�S���%˂�닌���pO�_L8H�f��܂�̘�.�cS��G�z��1�hˋ���
p��R��~�;jn��Q�ކ���e�x��+�Ǡ���f@C�Q=�r{��j����Cd�P�8Zj�(`Dr�}U��~���J������ő8�9��w��B�'
b%�B��ɟt=}ͳ��.��̼9' P�4	�3�*�y���3uoG�)�j�8Ң%4p��4�Y��4z���Q;\���;��k��E���?U*qQ�|XR���N� _�*-�o�1�o�親xeQf�mu��cZ���BM��J��l�c��*�  ew;��5�[u��A������1:�,a�=����Q?z~U����.�G����B+�ng�gJc4������:"�6�wg�c��:�q�c�B5z5�����K�$�ǚ*�%`a���b��}&����N哻�\	:�^�bV̘��J���؉�$�i/�����+p^���)�v��C΄M#�	8�8�,��p@_��"m�t\�u�kTE�<���=uY��VVD�iQ�ŉ��ʯ���[����o���-���c�WK�𞑋��w�oŎ̔���XGEA�eφ���i��@�E��C!�E��S��V~��\a^?��B�{a�i��fe-ɧP�qp4({園iF�^F;}�z���
����9o� �v���[�Ƥ����z<�G�.B���PRAJ�aQ���R��0�.ʡ꾴f��?��Y�YȺe@%N�}/��g�&710���AB�5{�A�j�΀i�Q�њ�C8J�jf�;�&��R�sB��K��H���ll�]T��P_��Z����l����>�r3 �ݩ*���I��/�,C�9�6ޕ�hG�z��F�+��t������`eE^(��&�(Wڬ˷|sv�b'���<[�+��0o̗�4�hɾ�n>�~�!�6;Hg�*o��]ْ"�}͆Go寕!=F�i���3pF�V���u+�}%��H�^i? PpӠ�ؑ�̊7@�u�cLُ^[IxS�v5]JRŭΓ�X��@�{T�\Z�a���$p�3��ڣ-�N��W7�!�yI;C����x1���,���n��U�w�E��cxpI�ʊ�D�YAv�f3�񡓨G���d��5�W@/������6F�{+���qk��O���vȈY1Qᢵ�җ�#UY�(d�ou	��&�9�K���[urɁ86�z����q�����]�(�De�O��H ����m��(�DzEx�������Y��|k}g��ZiZWw���H8�n����>�
�8�{�7|^��]��&ZK6�_�I_'�e���l;9Z��q�q;�х��*�ƚql/[�����K������i����Vau��iŰ�_��\ݎ�
��X����Tj{��I��̱�	��25,r��w�`F� ��M�x&�^=���� �j�A;�����dY�JO�ª~(��6r��!�M>���b���;
�����s����}�l�j-q�@���|>R8[��\m;�k�3�Q`�:dƾ�/x����k���������?��Ɵ��_�,x}�.>����Oڏ\�fW`�33;��AJp
��,��n�G�i++ޝZ8* uh<�[��"R� J�o�K�?�/X]����!J��p�x�m:����і��1�1� gh�`��?	u�of��L˓��$���$K�Ÿ��yOA�(�1+�TZ
a�n���1j~�1=�9�m���B���WiY�/YE�#k�6�O���T,h���A��ES����{GT;W�m7W)3�^T�`�l�D.s��g���px�/��E�n�&�'iף�2`)�O� ؐ�*0�9�e�B�и<�3���V�b�E8�]��
��8�X�DX�eLcQ.7wz�M�=1��W�/��Ď�xA�Z��FG�Dճ
Z�ޒg�+�{b:��*s�Y�c@Tʄ�0�(Ԫ� �G���JL�9�!�h��m�=��2jȟ�]g����C2�w�.^"x�{�p�nw/�C�h;�vD۸��i�ydr?�`�C�]��3���0�����
���/�Y[Y����&WLO f�=����������J�i�M&y~��s��7�i�pF㿪��Ƿ�����P�^nAJwX��ڧt��RWjp��N1�[�'��玂_��!�ҿ�8�B��h��p�.�W�9C&L���߅�c�dV �y���s����c(����|��N���	�L� ;��ށ�24�Q*�_~v�s�k0F�|�L휫LfG��������&]߷ŋ�}�sϚ��B�g����˭�S�����
_Yhg�u��\���C�«7��W�?�H��*3V?�[oOFk��@g6��.wV�X�3�<�Z_��ɝ2w=S�>�Ei���C";1��d � ��!��'�%-"MQ����B����I�3�7R�G�����~^a�G<��.z�dʺ�x)��(A�e�˂[�'���R;0'K@Q0Ž��L�c�r�1�}�[hx���8éA ��6H(�����+��c3��3^u�;*���%PR�P]}o��̤oI��e#h4V�;G�v'<k4!Z�Z�Q�Z3z���ig���m!��[�~�sr�hHN9�ب�W�7��à��(|m�)�ȝ�DQg	aSw�	< "_Vi`��w(�UM,?@���Eb�>0"�`���OO�<%=^ �rFԞ��dMȊ�yv,9�d�7��ـ��؈�%���ԈO���yP��G-N*Ê��,���&Q�[��V�oA�H~X�s�NĹ�~:��k]k�/1A��	jae3�����!���0h����V�V��0���;j"�t ��3���Ī��7���|���f��~f�q�O�n?��w�\p�$_9�}���Z�%�F`��t�r�'튘t��8��ȋP�=��A�v��c���$�M4���Z��ХE����������&(P�LV�D�S����ϛ��3Va-�����({C�`�%���Sğ��^Tk&!����� 5��P��ݜt&���J��o,�yJD�(���zxہp��S���%���$ᆢ��Nq����Mh:��i��p��c��ևQ�G#�"�ug��꾋����m\Ӡ���^Ç%����HL�Mr��\�L/`�s��&��N{�	��9[ͦ ŵ��2�I ����荰�98K"KW!����䎰���Pvl��U�����{�m�X��Ӳv�L��'c��|C��D�j�h ��X�4��m�$���~��nܛ������ |�� ����q�g�5q�1J#��zY+�in�<�U�߇�X�������տ�,�$"����uz9ˀ�EjTbq��B6�:Sg�Q����}��=�F$�b���E_�s�c�0����Xz��O?�L��j-k舛������U��05Z@��a`iB;m��N��U��%��lb�(�j�Ǧ�W�����4���s���w�N��w���i�����e<�i�7ѧ �ˠfH7��ޓ$P����R�V6��/�i����Ky��;�N�($0�>��	<3���L)��3$g�3��~��K��]%+�b��z��0V'"�6f�@�p�`i7�'��U���a�T^�Q3�-j��x���H��J�����<�����3��Y�&�����\Q�������.�Pf��S�W�he�"�Y���S8A�6Z�nD�P����=X�ɡ�sܚ�YxoaW!�S����	�G\�H[zY��N�
]ԯ.�%�:��0ͽ�����׀�+� q�c��қ~�J�%R�*VaGʀbt���=��4	H������*v���L݊m��5oJ��F�Ut�3-�8
6[7=u
֟=v�������B���e��!N�8��=b�gg͊��wE�7y䛯���y;^ņ� D�6\9�$H8e�c��B99O�8�X�냪{����X�ʔ`X2Uxh���C��ᙕ����A�3�ɷ��6�K��݂��C��pL���߲����&��y��#WW�}�h�@1�Hȉ���\� ]K��E�W�	�)7�fOkYn��+&���/>4i��(�X�^�8�������m�1,煌{�b���5Nf ��������^=��͑�㮼\�%��t�L6����P�<��ʾz�zZ�NL�KU�^�4�4v@���dAfhK�cS)���/��ؿ�<>�
��M �_:ê��0��S�a�0�B�G
@#ι���pf�]���G$���>�iIUV*�y�w�&fZJt��x���!I��)�߂z���FCD�nj�^�� �drC5���o)���:+FRf��L�Z ů���N�W�
$��r�� �$��YI���Z��D��S1q�Q]�_�e�K2�M��ڥ��-ղh@�Ew�H�#�Mi��
��߭W�I�V���������j�|�A�*���R8,�@��)��1�c�!א|ީ�?�M��矼?��4�2,K���EG�E��sꚲ��)�"t#�����q�L�'��Ʀ)mg���?�����Pr:�ٖ\�*�.� ��mA_&[��>��ޙxI��ok���+�ɁY1 ���q3�e����m7��ړ��c�-�������[�+8���(R�:���8^� ;�/�C�X��_5��乼=��u��F@v�b��	&&�@��	9hn����"_Ȳuj�9'�{Knp`�tm.�XɺT���z��	��ݨ��Z�t~��O��bݹ+�5tY��^ہ8a�����7)�7�:N��6���e!�������>09�'y;��j�Q )�3�T��#�sU�Q>9�6�>��05�8g����C��k��\w�A�@v_s���@O��'��)��P?�hFճ9����"�:�Q��(ڥV���w	e�t9�ْ�u"�D��^�Ǆ@�ǠV���9F�v/�I5_X���%�u��i�
�^.�m�֠Mk8TK-<k؛�u�?O�p1(���o`d��V�X$�Fç�31���$��P��$�s�&����	pE7�
�5�&�<�A�"�f��f�]��z����z_0ѷD����~g��X�^Z({��K���N������w�|���(�L�G6��H֯ys����@e�>}�O�e��LL�� �>���w2�d6��c/ ֻ�}ȡ�Vـ�~��B;�ͦ�?�OCG{s�(��l��^زN��_�`�r�^/�L�KG.�|JB6)H4�s��?�������Ț�O�����M�l!o�5��<P���.�˔;���--���2�fd�,�K9��T.�Œ�$�B�y�5���7C��~uu��uu&��;FY�_��k���H_З	h52�o��>I�� mV��Z"j��I�%��i*���e�y�@���2��0Y��ŅM�������G}�+�?����r)/�x�#2�x(VٱF�fUz�/~X�kMV=��z3^����[�ֹ9aK���ĕ,�t���Ǳ�tO��JoI�A�X�Vޮ�]�*$�"'D����p�	�GT�a"G�;r=�8�����}4MC����>����7�Ch�P'[��r�fv���!^��6��ț��>"���S��m/b�3ǉ�̤���Sf��Pi� 7����D{�Z|h�E4��aĕ����)+��Uo`�-��u�=vn���pb�gCL@�����Z6���<8{Q�������ʮ7cم�*��~�M;JC��A���Y�[c�O�|(��>���%<9�H"y`i.6���/6�8���Ct����>`	�xT�*H-�I���3:~��0���_e��ͪ�숳?\¬+�X������A�:���{�Ģ����ܦ�᜼y��݁�<(C<�x~i�b䤚�h�/�A5��sŁޕe&�ƿ�Q_�Q�[�|�>����&�r��(����BY�,�S�4���,H;��y_5�	�������^�?H�~t��t��G��p�@�c|�Vn,>��Wz�:ɣ��u#Wm���p�{�s��DW���t����ҝ�')<"8�����W�Cr��\Ƥ�-��uS5]����{.i&��	X?���~��N�:>F���ۣ�t�t����FMS�O�be��$_�Q��e)T��R�v�U�z�y�u�hݕ�e��j�mF:�4g�T����g��E��$�S�9�^q�N[����V�ZڞBu�\���*�������>��>��+^΂�/T���N�{,.�s�YI������;�$Z���B�'h!���Bl=6[%�i43~���]t�Q���H��X�b3��\����xv�H�j�HZ|���y)�>}ǆ/�������d�N�	G���;��2O�"�L7��|����d��H��J<�4mA��ypi��J9,�5�I���E��ڜE�""q��U�Š�lqK�o���p~�זEĻ�M����Q*U�錌FǓY�>m��0���1S%��獛������6@v��!3�X�q�T�xL Z���(%� x�}l*���fsj�x���uԂ�TdS���}�cFi����|^�{�!{	~L5�_���|�sz�+�'8����HdWܱ�Ь�/�0�ʩW��*��n�%��Lt�Ʀ����W1���#x��Z��ְ;eq¿�8�nk?�V�0����-�j�Li���ԙ.�o}��	�N�c`����:��j��+sՑ�s�p�׌=��]�h��YW��	eԇo�trJ�L�'g���B�����Ipm��_�u�%KF��̰�j��xy��bn!̳��ṯ�$�#{��~J{%��c#��n�DZ���ޥ��ws���!�'���ϻn���=-�����xhL �?�$��������Ԩ�x��˄~��X@�IU�������ܗR�l�"������@�����I�)�.֗6V�b�{� ��%=3b��ݱ	���t�u�Z���iJϛnC��4
u�{'o�3&� g���c�ev�^���/�s��c��&bu�.��ҏ��!�ѪFP�B�JY� S��'��Ǒf�`�b9�fjez�-$ɥ%jrUH|"���ۡ��;��H6��l!:�~�m���1w�P�%�L�Ck<�?�ų��Q�+��İ>�k�*\m�#�Z�A�n��6�y����06�hɬ}Ǭ����=��ad>�|saJE����d����9��
�}ݘ_᫔֜��>Lt5�*���
sN�P(�;������+6y
��a$���\E�{��S-���5�\�}��&�O;B�0b_x�_�S�Ei덯	�R���1���*�m*ل�j�{��Uo�&ԗ Ё��W~Ŝ�����k��C�A�#ޣ����'�ڀ���+�X�\�������-���?���I���q3�;󩑾��G
X��d��2v�yh��j��p|t����\	��xt�T1v%CBEZ1�%�-Seh��M����=d.Qn#iG<���uL4�r�Y��/J3��|vb�+<UJe݈}3ɩ�f�g��-kh�ja��C�,�JC��XLMJ�*\!$�e[m*���M���PQ���D��P�����#nj�Y��!V/��/��j�-�i%�g&�!��%b���oV;5vY�b!)py��|�z*F�Y��9�a�\�"20�veC��J��ں�����FRS8Ᾱ��rq;h��c6�t�O(6PIL�z��x���h:q�=�=�"�f�E�#���ޟ�B���܌윹�]]>���x^ޓC�����6��^�6��x����������+.��1�M.��'��Z:��lK�#&z���lOva��>L̡�q������yz���w�dF��c2i!��)�O�l���&�R���&�"E����@�g]�^��<�r2�x�:W.�Vƽ�+ Y��i���WFo�R�Ͼ~�yoDP�n	,�W<_���2�k_�i� 3���J��5&��E���?�A���*�������4}s$�;��ܑ��Ͷ�Re3�A�s'Es�nx:#���3�s_��'{fv�Q�8��m�[`��
y����1q���x��s���p��o���ݖ��|q9�;4|��"���cJN1�G��*�~G�8�"�`˰��" х���
�˃[����r0��P�ы���`.c:0pmQwj��qE�C�%���c��G�S�U�`��� 溈�*p�/0�U������|����y�Z�٫L5�eej`O^���=I�}^`� '��j�j������l,�α��A�0���^�^y��J�7@n�j��|僔ى��H|�*E�^�4���m_6,�B)�);�d��"^@ƈuS�0�n�+�M�TlkĭAB�Z�\{�g���cn�|NW���'`�U���<XgtM,(���I���Bub���yX�����m�p{�"�s�B]�̛��&���[i�P�Y�lt-��JT���
4�[;� ��.�L��!���ڨ� T�x�5���g���x���/`��;8�Jn`�?`[e^��[$��n�
4��x�p��D�Ԡ��օ�zɺ?S�S�N̋�r�]�0�吀̧]�O���aԾ4��9u�xi��o[~�V�2�"Js�H��(e��h7}����x���K���l4p,��]�˒�!��"^���M����ԯ�ޅ��)�ɭ�%cmL[���<�� �j3=7C�r��_m˸B��^���<�in��H���I��%�`�5�1yb<��G�"�\���)��o)�UA�H��:E�Ľ�b41i/.	�B9��+����y�_}t���UO�[��m��'r"��D�U��4%{��[��H\r�����Rm4�j�Aς��jr���B�L\�kjp��'ثi���Nd艡��bL��H�Q,y���N�__��6q=W�=)ΡcJ=��5��P=ʗ����
FA9����Ԅ�sW�#j��5E�5^b3�m�y�i� ���6P!�S
=��ē�)��I�T����]9&k���̂�=
���@�>Jb['\���Gr����"a�<�.�I��>q(Z�e�� ��ӈeػ�����C�3�F3��"��僆};^BL�Wɸ����
�������!ø��b��-�� ��A��4]��@�{����~���:��Q���3�uV�-���kG�L�bG�;;6�"�YLR�;���_�գ��f8^$"L��5�}��9M��W��c�&�otp"b����!����GpM_96��97�q�t�c�\�Fr�"�w�4 z�\SZ|݂M޴ 9 )1�ab��Ļm� d[�^�w7���@Ĳ�9�@�s�m��6i�%�=M��$�&y��?K�*��DE/<��b��I4�7'��JT$�="p��,���$1	c΀������.m;��2���A�=ի�vz�Ls�Tfh��|��ޅ�=�k�`^�-�x�hx�?�/,2�ʼ�V�0+1AOt���y�&�����ˉ�'X;:���#�hn���D''h����;	�^1��M}ӏL?P����13ꘅ!��S���_g:�|�e�S��s��b�C�MqK��E9�IT ؄�b��r��.ՍM��+�W�s�
��>��p����U�[v��@���cQ��:��-��q�?���5?�i�״�l [z�8>b5�Yo��U�-�k<����{��_ܩy�=9a"���cc���%p��ds`I"�n��������*+@3b�p��K_�ӑ�e�ЏRI/"�5|���{<n/J�m�u���w�J�fgڽ6��a������9p�E���a��Ù���(��4�S�R�s�rZ�N��7w��3��w��+��K���)��~�i��{lo�4z�
�]�*ƽ�)��@��;�q��J�0�?H�]�7O��[ oZh��t{�WFш�O"S8#���8M���k���o��Y�'�t���x���2�i�"\�Zǭ�)Q�K����/L�X��A ��>���'����Y�<�sM�b�j����H��7JxX�)�i{�{�p��DGϤ@�q��HM��-�9.THF,:j��:�m[5��ݵs$Põ�?S�:B?N�	Ejb���������Y{2�����n��������N�G�ɶvΝs�A*ܴᖑQ<㔆�� �r�$ɳ����G˴L�r�޲���=$�=�;�6q ���謹�����jJ�C�X�r���$eR��*fϝlD|U�'Yƶ�a�t��	�o|Lc�X����D�y�[�{���δ%n�A�pQ1ת|��_r��Q	_��]+J�8^w���d����
�0���ҺY��`fzڴGn%m����s橈��/���O{ln{���,������fp��0@�����P�Y���+'��e@�� T���c�I�5<5����riΤ.4�u��s�L��z9V��SP��P�Dn)����8�~y�i���i�;֓��yD$m�h��c�KJ��yzJ�br�z�ԅ�!�P��Sb�e���q�{���	��H�P�A=3�@������cbe�s��<��-�ب��ZJ��I<:��,����=��5�D�ب�_��`џɜL!�ng��(he���T���]�3pl܀�By�ǹ!���Ë�T�"������|����m�D����p�_�����:�u���Q��0����[NC �+��ĂZ�Q�?7�.�JJy`),�hj�:?Ɍ�n�O�h]��%�������ɬ�>�C�Y��$��ʰ+�;���.ܬ�-}�4V���Ƌ4�	��'oKw/�X`�k�F�8�7M�Y�N���X���S�����W'#��+U��V����f��h�T8��G�2{���2�Rƚsд�n�����D���{t�K��TS}KX0��k���@<�o��1��c�6���u��/rtu�!㚖������BJN���?D�ш$G;��801d`�5Hd2[>�@��i��vG���y�����6�w�%��$
w�*P��mܳuT��a�>9��������7ȗ�����?IpbZ�=zO�U�\E���(�暒�H�a�r\�d��8��\�&My��hu�U�0:�)Y�ݽL�MSߖ��Gp�Tˣ�I��m���,29�8��ڢ�`� Z�	:N���p���9wJ��V��#�`*��y{�~n����E�Q��t�	m!{"��Vi-/V�U��9��"t��dG�H���gK�5^uS*�ᔽFq�3N1� ��C<��(9c���كL@�A��n����Ao3`T}Bzw��sd0?�1�����u ,���"F=1�5�ޫ�ds������UK��=��"���Oƹ�l�7�P�8�ǿ�<��5�6έ�mpw���5�P:��Tz֝��3ß�h=U�r/澩D�#	�O���r<��P�g5���O��2�:P�F�݆"���<�H��1z�ƚ8�z"��dbEp�5�p.Hx�Ŏ���+��(�ezzd����O��� �^ǐ��}Ӷd�U�� b-��K�>��?��(�[��N�e����16�-����R��yl�%��^_�L��N	]�L����<�.���ǜ[�w��Ӳp��9�.%>ٯ/�'cɝ)��$��P�0^<g�-��F�)�3����;�?0s�.�:�bD���䃢g��^�M����9������e�nz�^JM�$��[��ǹ�:Өt|=@Bs�~	+/ѠK��-��#\({}�f��	�av��ш���e[Y��B�t^n^L��8�:;I���l����*#���Z��(��i��z?6DQ�$Z��
p�)�@����~��O��~�����}a�0�<�}�`�����u˄	���4YI��f�~V$W��r�
3/u.ޕ�ȣ��� ��܅(����X2c������%�J'3џ���X����\�(�-�e(�;�S�~�xљ�e��jM���#� ����!�z�Mmt4���������<{]^���"����Q�S*I�*Svl�ZZZԞꂁ�,66���=\�j#~�-Q�Bu*؍�x�0*N�G;��Ad>�?�����.����rN�e�V338�)p��@EU{���y/����4H��C�SوL��	��}F����<c��� l��㐊x�T`���5Cl�Iя�u�x�t�7Ҙ.�d��� ɷ��1�'ae�z�����l��tZe�󌚮����t)�*�ef�	w!D?�K�R]?l:�d>���H�#w+sI.6ł��&�K+z�i8p�Lt7\C�	@�������([mH��8�[Y�C-3H��=B
��W�83&� |�5�n%��-m���l���+������?�cq��S=��j���P��k����ZLd�/�"=\��Ԭ\!��lD��;.�}j�9��ֻ�՝@5 ��6�͑�UZ�˄4���:v�k��kqo ����		�c�m)a�����`Ԯ���Ȝ�n��k��!\�	oP����Y�Š۫�S�g�,4�+��K����Sm��9�\z@!qq����XDu�n��/��^��B� ���zM�%;v](�+sSɠ����\��&��='T��I�"Z�ڜX�c��T�=x�o��
���!He���\�T�#�e��f����:HbR}	kO�nA�t�y�D�b*���U��k�gҮ%���glM�X�@���ݧ�W��±qC��H{ �4[`Ϭc�(��8�Q�}��%��_n��<�r�(B��j����:'Β��Ń�pKq���Ǡ^M�m@^���?`5�r��3t?T�nTZPG��Q���"�a���������E	�iJ��!���?��}'aG��_-��vy�.Io�p�S#���S�k����CO5w�HtK�
��R;�P[�|!���{�aӂ75<#�z1'_�B/@x3�βiB�N_.���7��v;�`	�\��D���FC��p�c����̔��S�h��x�3�J�����_Zc�AYU��4��Q�25�z��t��¼�y78�+���*��]�Y��#��Eǵ�1���?0��(����p)5rz��Dv�g>�N]�MC���~,t�N���Qo��C��jy:������X���f�(|�Z��6��xhl���-b��A�p��F��t���ёn`�jU�uʎb���~�R�����(WI{��W���"�n�GlNee; �x�ہ�jq���EcЪj ?�&��Ry� �;� ����}Ϙ����G^ŀa~����=K�����ʿ��)�%��zϨ*�$�rڇ2R��wG��ƣ�+�R��^x��	���L��
8{t�G��0�K�4��$�`j쎔TJ#)���2K����±5c��}�+"�CxY*�:�?4�4j]�����8Z���!��|����^�F_>�R��(��X%``/@݃)>�Ԯc�K`"�Au����<��Y���z�� ]pC����c�.��� :�U� x9��^�/���[ܧ�}l�����L�Hv�@��K���i j�?kg�.�@���%R��?�����I��&���]�+���d����V�����́��yI��o�S�Pp��4D��Yo��3��;H��?�?���J�ꜣඩF������2=��*��l���B�8�+ĺ_�J���8�{q���N��lo'����+y�5|��*��f=��B,&c�Ge���36��	U��	�b�M1ڠj�{�g��V�����+�����=A�\6JR8I�b__����Ӊ��~��ڙw�hBo�/��[�/܆�`%R0 ��si�뻈:x��ZŻ��[9���}NzfagE�-F8W�����A�����ֻ�
e�}�~X.H��x�<˧����G�]���貚�t>]��n�����
$!��~�O�\����r cӛ�@��@�l��:��>6��%}��� ��M$���+�4#~恸�.OB�{���d�ӻd�A�!2�Yh�G�^z��ݙ>��A.���֕���(�"�de�^k-V��aS|���]I����<'�#�g݉�p%�Tx�����ȁ���xr-"7� 5~&��?���4��~b� D�EZ�h�Y�F⼶'�2���� W((-��A�Q/�n`�\��V���d���q)��T���f�����9�M<���.HS�{��p�q%��s���%7�x@t�b�r@q8�f�u2��;� f���	��G�p6���	3�s`�����^�y�~���u�&"�(��1�ŏ�.ڕ�F���}ktݴ
�`�sq�(C�U��ŏm�\>�_Kŧ�|�d�����U�̈́��~�'���{���E:3������\�U��A��ؙN�Z�4��^�������t��>��O��o���ݧ�h�YL��*��YsIp��uG�H��C���ވ���[|�:A�t�U��,�&T��Q4i��[A0����X�:D�K�O�t���wO��#�	�)�㦁B]���_~�
��0-WO{O{./�2<|�e�KP5l��ĸH�����11��U��u}���I��C�]��{i�u��m��|kU�[S5Q�d��e�C���(80�Ͷ�P�����r�ɯB�1ߋd�� ��1�⇕].~���pl����������f����83���o���� w�{��J����/�,¦!��Ov�3K�VI]��~+�Jb�v�~?X���e��Bjj���ɇ�e4lL+����V�`%zKf<�h2�7kϺg�6�K��3	��0&�'�s�GhX�����B{7H�MH��$��U��N�(��q_�+��6�(,!�6��(���U4��/��>��N�a�$�vS-��=uH��� �\#�Ѓ�1#�u�cM��9�ó��2̾&=�H J�I?v<���f����i�9r �;�k�oug��b{��6����C̼�rYj3�N�b�\��]���Oܗ��]Ѯ�I4���D�.�|��%T#͐n��st������2#�>�C�#�����@g����ԃ1����&t���8Xޫ��d��l���&қ�I�����.�<e�ؐ���Z'U���fa���N�	 nr3�ü`]��X�i�5��:�V����g�lq�����	����՜K�t���Q�����WH�j."�@�j�
F��od�j��ı�0\J&pEqO��Ȯ�׏���De1�������p�S����&�z�37[tH	
�XْM}g�'�y�QzI�v�qZ�61�7h�L�rr���Ǉ�[��-�I'V9n��x�øg�'��Y�Y��=���l!�2b����ǩ��GL����9�g��|ך��l���K~ 0ش����zi��/����i5K�<�AV����~aǁ��3��4jW�"����� �v�q�vHnvw���}���!�V8��\h�$�)��7��.�(%,!�X�쵥��5c0��;b�c�~�WR?;ʈ(�<b��'i�S"-������Hd=E��Ԣ ���R\V���R��.z3��eq���m�GA ���%*Ky�D��:�����}/�;0J�0�y�2q_�p��N"�|�5�
]I�"*�L0�}i�f��ڲu|�Oeu�ipO�ADL�{���O��x��ó��f)!ra���Ҹ'/�
$��`�Cp.���1�)_f~�~'}���ӆ~9�0ǭ �v�b��ViL���u<Ո2r�c8�bJ��Y�\�|���	��t'mA9^m
����m�6���5�k�\�<�d�ԙ.�"E� ��ҹ�`i�3�WHR�K�ɺ�g���[��'q�����B6#���Sc�0P��}�̋5�U��vפ)l
<�b���3�Ε��юmz;�u��t�+�9h-���/���\A��X��!��_�MJ���Ҷ�҄n�Rp��ϊl�O�\�M��y�>u"���*bq�%Gǵ�������p}�>g�U���y���p5��3>$����'+��;���%�8��s���g"Z��/L�~
�^���o�o���
��o�E�!��hu�Q,�B�S�9�=r������BY��r2�N�?%�0%�֯��I�*�1�%a�]��
���I��`8����=E�eU1������\S]C�W�)Q{��V>j�Ҭx�~6����,�G��{<��1��:k��v���R��?�@���=�Z!)^�C����ô9)���췔��x�;���jJ�t� �U���נb��I�śY0��;����X˪/��e3�4�����+טq�3�!ė��@�>3�<)�5&��f2lġ��E]���8��Gqp�y�{0��k���L�������Kq��o(�>ݘ�,Tu�c���<G���ҍ�s�?D��9��TҢߘK:�����H%ߞ�^6�A�d�C�t�
�~�Ċ���_t2��
�i���aL��1l���:���yP�$����؊j�0;r*��*�ٱ5��:���cnzT�N��GU!��EP��#"S��ї�{�|����$D�ё��[�vpT$����0|ZX�ן++��_�x���>f( ���7�t�l{AKqjf�����ۑS�k�o�U�ǼA��Q���K��\����%��� vA���4�h�2�7����(=*F�8~W�Z�B��?D�vO6�ф����Ksr`���1v��bZ�;/O�y|�4�eA�>�vOW��T�`&ⱚ."�}�*4ұõ�MÖ��Pf)�]�@5�$Ž��R��=�T	����w !W00ϓxw��~U%��[#���0���Ņ]z2�(��i��{p�0��+��ֵ�Q+ʨ�d�~� J��^Y>>���`ߖJP�U4�jcB��p����'} G���9�/��U�\r����p\�m@���A;�HyGN&mόC�c� �MWWmR�2"���H5"O$b?��{̿]���W�Ic����u}�B:G,� �#���{�����nt��K:`ϸ�+k�(���h͹ΎN.�xt��8q1�YL��
�ty�U3ϩ@�d�������=
��Tg�d���R�f���k�����'��y�	�۰r%�U'���R8���H״�&0�b��M.�o:�̃�*M����@&���$�2"|��J@��˽�!#��ԝp��zSG�ob��`Ed�1j��d����������a��3-�K��$s��㥆�8 �H����:.�%Ĕ@�H�B�ڽ ͫ�pFt����Ǯ61�ZI��dIAʹ�A�p�>y�`.["�/B�`2���W��wts����5$C����B%Q(��_����K�E�մ��������@���u�C�匒�s@�����~�?MW�Z�<U��:�o"f�,'�c�>|K<��V���;Xl����t��g�EXP�.ւ�pn�yc�R��䗫>�6�S�Z?���\����BG_�{5]���ET���i���w�u��A˩P�z��rۑ�r$��	D�e�9W�7&��{�3���QB�1,��C�r�bcl�T��&Y{�=n:'��������Z�x&w��H�����l48���NP�����P蜁Uʠ��i{Z�B�ٱ���T(wơ�Tj�@�Ir�iP����H���;n>�9�����i���HH��-�X��!�&�RLk5C����q�w�"�D*h@۔��V�rx������=�ЀA�'5��%��N�����m��5V�����T��ғL��n���C���@�<�F�Fg(Fd�z�r"ڍ$X�xy$��}��ǷI���4�c�4��a��P��F�!���n��+HC����Y�\��Sd�8�[Yh,)VXT(1��p�O�-H�lw�}�:г�jJ�y����s��Ł���^(������V�h�$c@���m� ��E���ۭ3�A���EeQ��*0ڦl����q�i�f��Ls�{�`	s���`B�Ѧ��WC��d�Lx�P7Lq��v�n��T���� �k�׬�[jЊИ��
F������`!)P8S%N�j�h_�p���^��|p���|�f��� qOϕK'Y�4c7��LB�ph�1�V��7_;�9���h��)��ݱ��!�#�-��w*!2`�9�:�G�@�,���['A��SX�����=܅Ff�.��Փ�,���=�(`1���9#ۘ_�XjhS���.���%)�]\��-���J�C��}��ܘ�2_֒����}{�Rt��:��ׇ  }��v֌h?���S��ֿ�x����E�0x_(�9��w��n &�ܿA�v�αRV�l^�&TI��!N�7�X���'G`ֶP�ꑳ=���
�;���`p�fH�A>�V��R��v��T�Dyv�h�5'�{�LK�?ܛG�gL'����d��A e�8�u'�e�J6���'�-�A3��<ý�-�Y�y��|��g'�r�*-��$�w�%M�����IQ|:��� ���6��q�I�>٭���t���N�\���w��S�%���.mR@S3z

���t�bڜ��i�C�>W�3�R��N�ģ)��w�섚bA���:~�"�wr%�VK��7Lr�IW�S12�Ӂ��M��G}HH�㚁
�'³��xR`>ƃ���%)���ed�T%���[���6ٛF�w����]�5{t���ɡ1�P�2� ����W !7(yq,M#�$vT&v`If�֠ek�v�ݰrʌ2�77���{u�����#������F���,��t��;5�k=C`(8�ևɳ���?����)D#�0�Q{��N5^�:�����WMi�#N�\�-5h�7Jw,<��Q���g:��"�~��b�(lv���#B<�X�(��Y�^�xGzT�-djE�rW�.�R�*�$��^�6�2����M��H�0�_g���A؜�<��awU�?�8��E*����4Of v��,i���k�Z;Qmǜ�S�O(�xX����)trB�Ϫ�6JǁH��J��Z�yc 	cw+ZFg8�k���x�����שW�75�}9��7M�dG|b��cb_4��ٕ�D���{��y�?�ѵ0�b�#?�iux���༉Wz�}T8�, �>�N�%P�_�D���-���VK1��8i�����<����d�Ho�$�'�L'@�0[˯�ś<�	��𙖜[��Z���q�7YZC��qV�RƏ�!^�ĢwEj��̓�&n0�dL"�
���
�?h�RJ���"��sX���Ի�&ľAм����4"T���$��f&�t�\�S��6�}�ٲ	q�{�����r[�G�9R{K����X��fb�lE��v#�׏��Աcr�ΨҬ�.�a���l��7��\cB�[?��-0���_%��w�:b���/� ��,��Y�4��e���*��>�3Θ[��OfӐ�UЗUO�����^����jӅQ�K�%!0�8��ޅJ���-�h�T�v��ԥ4������wd�i�AN�r�0Iu� <S\�g��&`����Y����+�/��F��滖������y���<s�B��H�R���%�k]���SMx�Vu���[�E+�g���s��4gȼ,ŵ6�`P�7�uX�����F�S�W�ny�_�q;�H�p���?��UX���g�>GP���`x�e�Ѳ��;����k�dE�u��B� �fAkC��E�*%�7�c$1��� C���^��;�w(Gf��;�`ɂMfe�R��A�p���� ��*&��f:�:!)�r�U7���M�M�-�T��Jٳ�l�q&Ԝ�����h��R���kO�_���7��%q�,�]�h5��m>�-�/�L��ʫ$��yS��0���P���o�a��٪8<J�'�r�6@f&ȣ��{~M�ډO�Mw�uM �ۈ!*%mr!�8v;���$��L;�h8��(���NoΉ"�	ֲ*�Ǉ���-��Lz���O��TaK�y2j�5�9�Y��W7"2v.�V�}�!��p�]B䢱��G�dZq+q���Y�/ck#�����Z.�Z.��g�B}�
��qu����j���O����� N����'��B�I<��?F�x��*Ž��7d���M9�-И��в��~腴�A��t����i�}Y4���L�`�F��a��o��-R��2x�{����_��R}���Z�~�{����؞P��z���(A֡ B��BB�8ꐶQ�j�Ϟm(���lJ\naW��YW�]����~����E�%7��v�z���R�Bz�o�^���!S0C�@a|��r��w?�����̛�i�i�-Gd*������$#�Pu�7������w2���B��� X��oqv�1@f~C��D)���`*�Z�i����'�����t xV�K��U���g�<.��P
����n�MH��!��4�"�M����.�#_y��P���1}h��%���F������ؚ8�2Sg�;�c=��"? ��ѐ/K�O' E)�	��5�,��/۷!������3+j{��׻�ېP^'�fR�~��d��e3�����z�ш����$/ը�8ᒶ�ɧ�zϿ�rτ�:A#cq:s��8V�L���� ��!������%�h���B,		6\R;_m/�:�����F6���=�Ay
o��=aWN��L��=*����4C���$\Y?����e����G�n'���B�O����Wc�F1���9OK\�]�Aʢ-��,���2��Ze��}�eQ�f�ȋ����a�Y乳�.�p���4����y�6�u������������8� ���(n����/��ILݑ�,iN�@�=��C�aJǘm?���ൗo�)1����~�0�+pXvG"����"��q�Q5��~�0?���t2�Ҡ��}����Z-�X�0�8�����,^�YQ��9�&*D�aD�Yn���nOb�MHq�h���X�`���UK���xc_Z�(�"�e�{�I����3�Wf��N�������Q<Mǰ����HW~*�Km�P^p&i��(��n���z��hC�=Q�vDC�橩_�I˼���;��X���y�����T�M;��8P+��V��L*T�4rq&�>tL�qS�>�Wm���� H%hEǽ��_�#��-ט
m!���l�ɢ��/��3t(��)�����!W?�,��[Xպ�z�*l�_>;O�C
~�b
�.P�]�v˟j�;�� ��m�?��v9R
��U����z��IDK�u֕l6���{������HU�^�D���AQ+�"�w�g�]����l܄�ڒ��j�\�Y�;��
S���@�!^��Q�h:�sZE��Q�l� .���K���!'b��A���7��#:�f@�J�"��N�2��k�}'�(Xt	2ȅ18��7��Bc�l	Q�&�qD��~��ik�G<�U�Ǳ>t>���Z���]{2�6j�ڞ�������I�%��x&a!�}Q1w��g�0�,��4<�pi�f�y���	vN����Შ�ٚ��Ɋ7[�m����$YG�Tn�g��a`�C^~(Zk��%=����t��`��?� hl\�&e�|� 'èi��6+vB��\Ό1VЖ� $���	����Q�2���{�bː����Պ�W�DA�s���ې�I2R��f�����U_�4� $�������N�?N���oϑ� �ܝq����P���8�e٦�j���\�4��Xh�@u �ԥ���l�jd��[ezY*>Y�Ul��G��80p{�ua맒��!M����vgCj[ʣ��)���=b��N����k��f	�OP�=K�ؙĸ�ڥ��~�p��9կ��7d���[��;���:���L��u�e�I���pv�_���!Sob��7d���i톮x�t{�v4H�4��!['��p�#U.��{G���S�����A��>���(J&�+,�hM� ��ǪM6T_����fҞ7)~1�ID���	�I>�Vޚj�3��Bx�b� �f�:G�w�Ty��;8w��b~o�[�J鬞z�HS�a$���7�Q���=.��E`�ջ���&���\0K$�9La���NF��o���@@0����Z7��qZ�ְ��ϻ����lJ���e�K@j��)�"��8���5�4�C|G�N͈Q���~�t���.�i��-y��QS/��>��o�?�nѴS<�{��0�0�b����$>Nʽ�%�M���ܖ�QMj+�+�D�:7��az����vgZ=GPp>ls<�1$�x�&-�}�|7UQ�9N�`qE��=��'Eig�"-�_xT�hu�2�����iy���T�ka���Z�z�x��$�4�Q�syJT,9zG}�!�no<�K�����Jfzpa�ܦ#�m�"�|#uF�۰c�ITʻdӚ�"yG��j�`�-a��P����_ �U��Ƨ��Ķ_���K/�B����`�w���H&?�8�ZZc�*
��P�D�mJ����X2	��l�%�eF"�����D�8�|g��ý$�Y҉���w���)!*~�||hl �h�Y�UL��>ۧ�y�_�o�
+��|�.?!Z i�ѥH�={+o��o�K�C�x�Y�4��B���!��z��9� ^��$�[2쐜��H>Mq��|���v���i��D�2 ľ.�6����2��H �m�-��j84���"F���^ew�`����	4�[��	�L=JR�
h&��,�Yz�����eH����s�
��*���	ll4�p�� >5_�"�i�5�6|ͫ��B�U��8k�����(F�c�<��&�Yjo�DD�y�&7>y.!����!��[���uxjMt�:�� H���y1u�?~(�a�:�C���:&D��Yr-Еk�o��1�}ku�B�&<����
��l;>x������ч�}�=��:�� |�0����%}��2�3x�Jϙ.��n�!�
W�j5�fs�!���)�T�f���h�%�#w5>8��?`M�a��?K�[9w��ţ
R����jE�7V�\X9?��ĭ��sO>�ݲ$(ͪa�����t���q�������l�,�|�Gp��s���ޣW��%~<؍��>P1�<�;���ƒjo��Ɔ$Gv���vM�0�NK�W��Y�������g �f@���tF��Si1>M	e��!��v���$)�!x��΢��lM�JǨ;��-������:�]��sgE�eH5'�A�B�[�y�I,�g&�=�N��PfB����r7���t���R'`�W��A�4�<|H>d�d���R����#�����׽RoaCm��!�m;����6�W��MJ�����hH�Hz�k���H�X�	F^�3����P�(��W��0��KUϾ��X��o��E��2��g������7zE7�3�ϯ�����糣��P��p��Py��z|Q���N��+��,s����ñ�@��'�2�I(B��k*�ֽL�Ghd�j�n/���������㳰����8�������X�������s�c\�(�zaɚ�����g��c��fl�<zj��4��?e
`ʎ�I���c;��5��:�����l�����m|g�W�r56��"�?�bRQ�b���u�i`��_�Е��'<�M�[9��/�&T@!��?7���/B_D7�8�:LJ(-G%��)l%���gn��վ��]	),&�����P��Q\�k;���V�J�>��V'���u;��b�����a'�+�h��+��g��� 4P���J9L��޽>��\�����t^(�F�)�g��V:�^�訔�O�,H���%��fq"uh�$��$�AB�ν�6��B<�����|��l	*��0����~Ď��"���u1-�-��Ym#L A��a<x���,X��'Ѓc��ETI�ruwLl�?s�P��դ&��KZܽ�9u �������ǌ����in֝Y�x�A�dO��'�1�:"EIqD5Ԅ���O?}��u�'�&� :
-�y�!�����Y-��t�)��l��������<�B�����m���{X�/���K��$�d�f\�7K'JA�2���43|�����Άgn����;@�4�<K`�iF���M�����I���$QJ̟��5Í{�:�"9��wl�k[�z��Wd�x�����$���=�Jc5�;�_��T�dbB�{�d<�@<����� I�^�~���7��A�x�~ɚʭ����p��A����]���l��&��Yq衕��3ob�^��l~@	t����^�{R�5�R|�	,�w~���u��J���
�T��$�N�9_g�6��Y��T��˥9F=蔙�'�%�:K�$� ���k�_[�Kv~)��<7\T�	6��R�ND#�,�~�1D�m�:M-4��P������Yl&�(X���/#C[V���7���$��[zOХ��A�9�a�@h�i�ﯫ*I�>��z�U�[뷚�u?��g�9�#����NP;d	R�S��wt(�h�x�	 b�~��.�T�q |A����9��]=&�K�[kfؗzjct9�x����Vz7q���nȆz��mW�	St��,�@ E��'>��([��k�	0�S���Jʚ����r��0�)w��'u�~��Q&NwӞ����@��"v����=uh�/��$��f�#�f��P���Tcl爻��#��j�%.l��~v�*8%/-f�7k�:� �ʵ9���b&7�w�x�>[���\#�����9'� �bHMj�-�;A�?�!_ۼ�%gd�e(�$[�fOs���
7鈵TPW�ĵO�����苝z��iw�mC�O^�X<��7v�����r˜�hA4a���VF��0%����lN�B���%6ߨ��u�P����xZv�ȋ��;�1��5>Uc�v�<ljc�P�F/e���XM�H�4��S����˟�kzU�cS\`?>���N~(��V�gd*7����;�+�w�-��ꓜ!(��N��H>�^����D���/[�|H	fxGQ���K��j
$���Ï{ܼ�묈/ɿ�_�i���E�1��6�=X���x��������O�!��"	^�t�1�Zu$���x���$�Su���R�>�
ɤ^�VK�5VD#�NH#{�G�[�{2��|�������K2D�"�~�Z"���n���Q�!,97*�]�)�g�<�V�ǚM�ӿt��"gOkŇJ��7:#Dwy�o)�ً�͇�p�Vc�c̚hE7�&��"9wR* y����%ٗkv�	��d4�9�,l-�7�cz�<}`#�J|f�,Nq:Vj� K�)�S9�`j��3�Q �LEI#�J��������>
��t�0Q/d�"�ћ:�p٥��^,AX1�J	����P/E>]֛��SP	�+��/ep�q3�A0����yK��IMI0.��#Z����h�(��ۧ�C]�����V�N��Pѥ}��@3�:VxX�&M��#�����R��bz.�n���D�a���Z�z~��ׇv5�⏉��r=���(�����*�i��͟8�C�7spS#OfsQ>���V􋉶��r�6]����S�*�x���$ .��*n'c�r
*��D�Ƹ��}"H���=�b�E�a�f�gC��E��Տ�*�&��޴���u�N�@��pWO��D�0~���\�ܞVm=�f|׽��/&_'4���V�N�đu��EJ�窸3�ں/ս�i���kE�q��ozC�tN���c ʆu�<�t\����^xa �0�`����I��5ѫ	��Ħ�_JZq[R�N(��:��»2F�FQj~�E�U�,Jي�} ����j#�ւ��Wmb��_�p��̣�Ú�Gb�ɖ�&��_����u��)�;���G�f���/K}̚�lo��&�L_�D����P�STHmP�A�2[�ƣ=5)!)O���溡����!�BOr�1���g6���o{7Ӌ��ٴ�����xȨ�- ������ΐ+�����	��0HзI�K��%�����Ȋ؍l�C	g=�/�r�:d09�H��i3���޼���ך�²ܰ�������_;M(.S����;�Y~�$y�$:�rX���2����@�3y3N�l�) �eP�P����wI�M���$�f�2D��@15�V�SiD�,��-و�,���WG�Ϗ���d�Z`�O�K�/˅�Z���L�����/�MH:�6ڏ{ޠ ��/3O���"�ٟ2b�$�|/n>��,�:@)�b���J}�TGI�1�����NZ��~o�Xhv��!�\�8y"f�k�����Dy���C6D�"�U�קW���e'���A��)�:��%�7�Y]~�z�JT�g/xq�S�,P�|f�k~�=����8�\ɋ�ך��X%Y��H�����.�炭9]	���,����jKq�4v���,��%� �(J0����i��J��T����+�H��������:$(�`��f��<W�(�9���9\��0g�f��T	�g�Y߳�8CJ��K0� >�~���q�h�p�A%�:�h7�ϩ�ծJ?�0*`k���1�.�#��#;=@���A#��W(�n9oT���on���>t��ʨ�ڹN�����8d��eS�j�ד�_z2��d�nM���eN�+�E�p�n�d-<���5�_h湏�B2Q_��"K��v6y�7��/\*��E6�W�#��]3BK�.�o|�ؙ�&��1��~��?&��v_�<((�E�^�Ǩ2�C����?����.�jM����ä�
���8o]�y��w{}�-�]��Ò� �G'�`�Ռ[�!�ʤ�d}c��!r��Ԙ��Ж&�v��*���2��"�����kq�{�V��m��$����5��l,�x���yg��� ����-0"�;�D�e���)Hq_��]�n��o�mfG(��A���#���=jaDn]ǖ�f
;�c�@��0�Rr��$7�]�]�$�Q/��/t©�l�?>��&;u��ӄ	�*3�����8����g�vw �±cV�x� �y'&��O�'��	��R!{�eYܴc�v������r�(�U�_@=���E��%0�̀���Փ���֦�:������.≙qՉ�l?@�9:!&��{�U4�M�F�Nx´%���FP�l������Dͫ�PǇ-�$ ��L*cg����#R	�z�T<���Ly[駽>��g�3ˈ�N�vۧu�*�M�V��v�*B���ڧ���[r2��\���#�gSlbch�n}�I3�\ "��w{gz���I-<��2kv�Ƞ�ՠ��*H,�m���䷎�?�N�_��P���q���U�� f�w�3�H�Їx�jD��}��z6�zD�2��/����Hc��[�,��޷�8h�Of�][�]}ib���޺���4�~�8O�sDO�n��?��6��A ��� �������0y�� �>�&�e0���h51NU��|O<C���7�1 e��%Dqp�\���뫶P2c�<@?���WP���ݵ9���c�zu�;/-o�P�\���Aw7n�S��(y�d#�z�M����+]���.�(�����wF���=��|�Z��7�r�vu
�a�K��x��+N����Ұ��F�~���[|ɰ�Rr<����?�m;�h�E>�46�h
;�X@'��~��g�(��%(p��v$ �Ɵ�t�Y��x[ZO�R����N[�_x	Q��tc3ә[A��D�(�0���	�<�.���fa���t���C�nݹ�`�Ɠ� �Ҩ�K�
��P��F	G:_	��UP؞� %���t�/���H��n6^�9𣏒4O�;R�z�>��l���C�Kj7��۰�͢I��c����UV��D�t��jX4h+C�W������9��Mɇ��>�N�hl�լ4���Y���󨘏;ᜌ��)�^���]ѕ�����]G�������-<WL�fTT*h�B#AR-\b���R�˅Rp�X�Ex��E��Ǽf�8f�j��T�8�y�è�O����;S.D����#p61>XVv��?ab��Pd��BT��ZؙŞ��-�;��L���m9 �*	����^
�+��k�b5 �����T��#7�.�2j�2�w��7"<`�!>���?�ݫlb�o�n@N>�o2��-7��C�U.c�J��%7
�S�U[(� ��4��Ȼ��a��u�Q2��c���_?7zVև�}Z��.3��g�}�K���D�b�����u<�!�+Lӫ���^���%A�p��o�b���B��~���ٚ��aKu�a�Я˟I�����~Ubz�����#"�c=��$����O�w%���w���+�1]���s�|���B))��¸r��� 0�A`��w�:��r{�x�{���<^L+&CEA�m3=�=;^7#C�U��b��;�0gp+�b�6r"�����Q�K��yt��%�\Ն�Y���JLyy+��bo(�}�+sgW�*�W�E$�88�!�׶u� �t��h�Xj_A�l��� ���Zb'�Ic��<���yP�6D�F�A7�fNS2�K}�r2��4n��e�9m��+��|N������ћ̈́�wL�m�Y�z��z[�,:`�r�pj�U��n�6Ϻť2���o�E�~�Z�X���hz>��N �J����E��0/->����q�aS�j����N���Ԯw��I���l���Ƥ�\4���c:�7�}��u��Sϕ��ܯ9$vh�Th6���(��B���"���6RM�9��$�<��0*�� �G��0.|ٍ�f0Ah��'BҭzHK�r��7�b�Z�@E�J�W�k�Y�?�U�_�/�n 5�J��ntnE�3�q����CA�PkN�rL��#���n;���$P��D���dZ6k%�5bD�'߰��w$"5<fGi��D�'�y���(���o��L�T�[@���=�����>t�N��`%�X�v�
�jά@��vӸ�ȕ*9ΏQUX\s߼V���,.)U]�Cj"N���6�%�Z��(�Q6��;L4�Ki=-������o�e��0=��Υ*D��a�ƅ�u�r����WD��	�PdKǎ�ME�}�����\���
��f���J��������"]j�F����yu�9�Z�DO�y%���o�t�I_p�xM�ގi����i�'[�;��M)���^Ҵm3���6ugT.�c� ��(��?�~)��g�3�q!կ�j�1�_��SpԾ�>���<Ls��Q�,p����E�	lGKb�Fc1}��-EE����=�ˇ��ّ|�z�/�Ҝ�'�
1r����|p��:x�ə�Ej�TD.��9�s��@�H)�E#�[E�E_Ǆ�	��|�j� "i�9H���: L����Z�t6g��	���r }�7����,Y��8NvD��z��a��S��Qj�T/�W�z۫!��F(�(���s�^���,i���ت�x�3��q���3�M���=~ݮ�3oړ+�b�#�B��9u�Uj� �ѓB˞�v=j.X��81p�.�����0l�,9�7����+��.�~p��?$���7h�f�V�B4�e���A��At����,#���3V��p���5��q@��w5X:V/�̡h�btx�Г�vI�V�Q#����x�8����x�,1a;h��YP�yʏ�xh�}GQ0���cv��x��iT_�!&��V�2����OfJT(j&B��� S�9hą7l��	�0�t��\l�R}<O}�9o��{��d$���f��:�� 4�K(�kh6�FAN�(
���E9}����?��,�h�o�U4�V W?�BDl2���ⓣ�ݚ���a��LQ"H�VdT�A���0x�^H\1�Fؽ�7t���U�u�y�S��`�w�°i�
P�����y�˾�c�n�QRB��~+��u���&�m lW�-�#�������e�+@��|��Tڳ�Q4�YMxM��� rP�G�j�ҁ����x��7���⦤֤ۜ��V�b�/���V:R����(�&k+�gyZ�X��O琴�D����f���`�+C��a���4jPj'�W�䮠&���:��_��z!>\��o2�ޟGΈ�39�jǹ�GJ�zaY����zU]�ܩ����tJ���p~"�$VH*R��g�S;�?|L��R�`>�Zs����*�X��!!H�B�6�@G}��u��0&C����!��~��h踎x)���2�,��ѡE8T��v�z���9R�����[i��?��u�p��mN`fZI�1"ki�$��-���_c�D�.<�Hs��s-��N�o��'B�<eSJ]֮���!��r�*��g�|��u��B53�
�v�=^e`�٫���V��E5]X���Fٞ�iw�Z*�ɳ�7y๠�3��J�'N>b6*��d�V�hLGX K؁B�QLxIR��n�G�LB����=�6ˏ(n�Nc`@8>RƸu�I�Q�i�]���'�`�C�ec��&�u"�0}|�������$R~>�B��5��A�xc��Y���I��t&���r|D�Am�����o��,5i6�	���An���}�h���k�)?P��N�ۄ���D��=�޿�Mp��$�y`�w�{�����ȇ�k�H��n�� B��G7��Aj�E>vtsR�^.�+0X�i}m��u�;��A<>��?=q���^��48W�<t�����b�����fr� ������GY5JfW���NU�eL�͂ݖ;U>�:�dG���O�&)6��$�������v�S>s��'�+�����ʑ	�1���z0^-O������H�o�8�wm�DI��꒮D=r���'��m}����C��;p��~���D��6C:*���꬜ !�g�ݥ�)Q����t����[[���A���rP.?
�� �^�����O���v=��Wb�tg��u����B���s� �iJ�?M��!*|�{�)�DL�!�?��>8	�p����$x���;ϳ��Y�.�r��
�[Fo<F��d�b�o�j�t���?Y�K'�������N�cí��{��^�Xio+�I�r>���FtX��ή�D�ۻ��`2jض����JI�֙6��t�-��zq�P����AӲ5M.y���{����*jLC��fST�?�)�cr�ԖK���
���_����630Ė�����C?q�3�ij�zʢ���#�O2 �o�B�b�`� #��U=�I0��~z��A⍜z�j�Y7Z{��4��i���p�8ǒm���[�f��rU(�!�&�mAGx]d7�
l���I���7S����v��Z{M�M�]��;*?~�L9�N^�(|���;,lyW�w��'HyzyPSFS9���,�����"y�A��{z���/���������3�h�����X���cJ44%p$W�S��|7��>��<K1\�GZ���v<h�V�ֱI���ZP�Xe�_�̇Ć��K�_�iH��]����X��AxT\�3C��Af>�$�K*WRJ��XgI湫L���`��jU@��Xrʬt�����4��'6�;�%�R��:�����ד�ykʤ[�Z��W�z�F{����!����� ΢^��3��W����M��1�3R�<0������]Nv��F8�R���ʦ��}ݣa�`Y�'�	���
wD.���g<��������.�3��1A���n���c�����ߡKo|M�$�&?Q��W���F�G�pO�L����W0�:5��h8=�b%�hGob�Q�J��� \;|L�Eif��^Ko'�yi  ��d�^�8W����-a���6`��#l��~Հ1��xϚ�_��ϭ��h�u�����+"�M<�����(}w�uH�\��K~v�e0ݟ(�ME_�U�t�WZ�N)��<�4F.;�FH��L��b���9��2�x�w��B�Q7��#Ŧ�o�9�ԏ���_x����x
[%rE1�- 1ش׷�Q��k�r�-�떽�e�'}���V�+�(�l��$L�_�g�%q����hSAr�S�ꔑA�2b��ڌͽGo��<x�Ѷ��lF&�����|]:)F$���]J��߳i`<����;D��)B^��$���l���F�����1���	'��p�t��%My=&���X_K��A#o����g�#P���C��@���$ǌd�]m	I. <Ŧ,�lf� *��ʚUrfϣ���|9=����j�E�椋3�>-n*]��1�$eO�~?�rϔ�5x0�rZ31I��� ����m*�'�Q������?0���8F8���ʘ�>k!���E����7E}n�C�Z0�9���	�$#����q��nY�]Z��d��Pj�Q�V���63�VC]�
���qۭ_�ٛ��:���]��6�p����֢��@q�(�Y��y�)m膹05�u������{m*^�j������ilЩdL]�O-��ݨUj���{�4�?�wui��I�Z�}�f~h� �B�������)�$��.���7Q��A�x^B�g�]`���4އ�'�a�H��*��b�N̊gk�d�LX��.\��:jE�� n9*��:/���
�'T�:��Ĝ����u?f9]���넇�e6T��>^�r}m��,�3,�˔�Im�_����S6t�]��c$��Ό�u��_?蹥L||��6�>�΁֝�U:M�V�l�̷�<�[��H�a���!(�3�1��(�{��2:�t�6E;YH
ge��~$��X}�*�i�v�G�(�4�W��Y�auP�2�#8��A���&n�B��߶	�\A�wE�eY)F�DTͮ2��Ւ�i�l�QE��)�jm�U����j��MU۝�1@��h�j�惸Nn�]M�0:��S�W8�p�Cio�����Ilԓޕ����℄�;Hu�R�oU5�^�΂ǔ����|#�eB�b�b�H\���Rs��J�ܐa�����K�.���I[�i)��F�=r�f�%"[{�����u:��P�3��1�v�������˒�6����_c��5�!6QѶ}���tb�7G332֚.�<�	â���u�<p��H�oп��u8 �,Ҫ�O�/��"�c�'�,�u8o��dœ������oGf^�Q�"o��$Hh������ʆ����v��X��>���kϥ�Yl������WW�_���O|�@���K^󲘈j��w�*�f\ɞ]r1�Wi�W"�x��9�,�e�m�7$Hl}�Sӛ�V��Ng�^����Ф!p��]�2�����c�$��)�����,�/�XB��+f'��G�
Mdo��M�W�T׋���CY���2�N��
�b�IJ�hۂM��R���s�$K�t<N>'oU���W����U]e�6�g^O*)iX��%��i�=��T��ᅚMA[��f���/A����
��t�M鳐�t��>�Ȭ��L�qo�����:��l�����ߺ���W��:�^�����\����x�᱙i ���wty�V�t'~�pV�8���"������kz�פTW��`+��kR<\�5�j�h;S�{�b7T3��N�w�0!�5rq+�y��s6,{� ��D �,[�����S⧘{��I�����6L����ֶJ0c��	�A��!���HNɶe��K�������9��.��I� ��0��jH����pT�����I���)6�
����e�8�xv��}y�ӫ�XJy!�6��]JE#O��f�(�A��w����N���k��Umm�\QQ4�ǭ�X��$֋:��?�5�*��;�@C��{�!�ׇ��J(B�7р� 0��ՠ`��\ ��}��;6����B�,+�AJ���V�
�����+��qI3��� ���� ��x��y��13	�.�����sp�qU�!+�m.$[�=wV�F�\Ӯ�̧A��f��z��`���0�U��R�b-�"�"��R��k��*�IJ�bu�T\E$�Y��=��#E%��@���ѱO�z��E�8|�A��v�;���������@��+8|������Z�΍�kN���HQ�)&7�;ߣ+K᫸
�H:�A��/5�+z�ݹ��='7��g��$߅���QAyj�k��ǵ�����c��&��W����/g�n�,Պ(�ި�\�,��+�7D�A�ѹA�s8���3�Գgɦ��ݽ�]*+���KSH������������r�Y��(�5~<O~�Tw��qhC�Y�Q3K)�7]��0��	W:���(k�?"����<�����X�1g���km͈!��(_�8�����d�^=�H�����W�},�<Fŷ�I�`D��+�@e`^ZI�g���E>7�� �0C���C�\��1�<Đp9��A;n_h���h�����50�8E�H��p�^|bǵ���h3\�N��2�[�j��mtW�j��g�z�h����&��R����B��2�:����9��q�t1h��@n��C�<jjv�_��OX����8�s���ǷI��\ng>+C��	"���OA@�-ӎKW�(x���N��|)3�J�c�J��#a�����ex���	�C�����l)ۤ��{�#����w�r�J�Z��<��=ޚ<��̿*�=�F�D�.يA+��}��)}�J$��|yo:y�@�