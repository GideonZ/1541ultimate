-- nios_tester.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_tester is
	port (
		audio_in_data           : in  std_logic_vector(31 downto 0) := (others => '0'); --  audio_in.data
		audio_in_valid          : in  std_logic                     := '0';             --          .valid
		audio_in_ready          : out std_logic;                                        --          .ready
		audio_out_data          : out std_logic_vector(31 downto 0);                    -- audio_out.data
		audio_out_valid         : out std_logic;                                        --          .valid
		audio_out_ready         : in  std_logic                     := '0';             --          .ready
		dummy_export            : in  std_logic                     := '0';             --     dummy.export
		io_ack                  : in  std_logic                     := '0';             --        io.ack
		io_rdata                : in  std_logic_vector(7 downto 0)  := (others => '0'); --          .rdata
		io_read                 : out std_logic;                                        --          .read
		io_wdata                : out std_logic_vector(7 downto 0);                     --          .wdata
		io_write                : out std_logic;                                        --          .write
		io_address              : out std_logic_vector(19 downto 0);                    --          .address
		io_irq                  : in  std_logic                     := '0';             --          .irq
		io_u2p_ack              : in  std_logic                     := '0';             --    io_u2p.ack
		io_u2p_rdata            : in  std_logic_vector(7 downto 0)  := (others => '0'); --          .rdata
		io_u2p_read             : out std_logic;                                        --          .read
		io_u2p_wdata            : out std_logic_vector(7 downto 0);                     --          .wdata
		io_u2p_write            : out std_logic;                                        --          .write
		io_u2p_address          : out std_logic_vector(19 downto 0);                    --          .address
		io_u2p_irq              : in  std_logic                     := '0';             --          .irq
		jtag0_jtag_tck          : out std_logic;                                        --     jtag0.jtag_tck
		jtag0_jtag_tms          : out std_logic;                                        --          .jtag_tms
		jtag0_jtag_tdi          : out std_logic;                                        --          .jtag_tdi
		jtag0_jtag_tdo          : in  std_logic                     := '0';             --          .jtag_tdo
		jtag1_jtag_tck          : out std_logic;                                        --     jtag1.jtag_tck
		jtag1_jtag_tms          : out std_logic;                                        --          .jtag_tms
		jtag1_jtag_tdi          : out std_logic;                                        --          .jtag_tdi
		jtag1_jtag_tdo          : in  std_logic                     := '0';             --          .jtag_tdo
		jtag_in_data            : in  std_logic_vector(7 downto 0)  := (others => '0'); --   jtag_in.data
		jtag_in_valid           : in  std_logic                     := '0';             --          .valid
		jtag_in_ready           : out std_logic;                                        --          .ready
		mem_mem_req_address     : out std_logic_vector(25 downto 0);                    --       mem.mem_req_address
		mem_mem_req_byte_en     : out std_logic_vector(3 downto 0);                     --          .mem_req_byte_en
		mem_mem_req_read_writen : out std_logic;                                        --          .mem_req_read_writen
		mem_mem_req_request     : out std_logic;                                        --          .mem_req_request
		mem_mem_req_tag         : out std_logic_vector(7 downto 0);                     --          .mem_req_tag
		mem_mem_req_wdata       : out std_logic_vector(31 downto 0);                    --          .mem_req_wdata
		mem_mem_resp_dack_tag   : in  std_logic_vector(7 downto 0)  := (others => '0'); --          .mem_resp_dack_tag
		mem_mem_resp_data       : in  std_logic_vector(31 downto 0) := (others => '0'); --          .mem_resp_data
		mem_mem_resp_rack_tag   : in  std_logic_vector(7 downto 0)  := (others => '0'); --          .mem_resp_rack_tag
		pio_in_port             : in  std_logic_vector(31 downto 0) := (others => '0'); --       pio.in_port
		pio_out_port            : out std_logic_vector(31 downto 0);                    --          .out_port
		spi_MISO                : in  std_logic                     := '0';             --       spi.MISO
		spi_MOSI                : out std_logic;                                        --          .MOSI
		spi_SCLK                : out std_logic;                                        --          .SCLK
		spi_SS_n                : out std_logic;                                        --          .SS_n
		sys_clock_clk           : in  std_logic                     := '0';             -- sys_clock.clk
		sys_reset_reset_n       : in  std_logic                     := '0';             -- sys_reset.reset_n
		uart_rxd                : in  std_logic                     := '0';             --      uart.rxd
		uart_txd                : out std_logic;                                        --          .txd
		uart_cts_n              : in  std_logic                     := '0';             --          .cts_n
		uart_rts_n              : out std_logic                                         --          .rts_n
	);
end entity nios_tester;

architecture rtl of nios_tester is
	component nios_tester_audio_in_dma is
		port (
			mm_write_address             : out std_logic_vector(25 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(3 downto 0);                      -- byteenable
			mm_write_writedata           : out std_logic_vector(31 downto 0);                     -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_sink_data                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			st_sink_valid                : in  std_logic                      := 'X';             -- valid
			st_sink_ready                : out std_logic                                          -- ready
		);
	end component nios_tester_audio_in_dma;

	component nios_tester_audio_out_dma is
		port (
			mm_read_address              : out std_logic_vector(25 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			mm_read_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_source_data               : out std_logic_vector(31 downto 0);                     -- data
			st_source_valid              : out std_logic;                                         -- valid
			st_source_ready              : in  std_logic                      := 'X'              -- ready
		);
	end component nios_tester_audio_out_dma;

	component avalon_to_mem32_bridge is
		generic (
			g_tag : std_logic_vector(7 downto 0) := "01011011"
		);
		port (
			reset               : in  std_logic                     := 'X';             -- reset
			avs_read            : in  std_logic                     := 'X';             -- read
			avs_write           : in  std_logic                     := 'X';             -- write
			avs_address         : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			avs_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_waitrequest     : out std_logic;                                        -- waitrequest
			avs_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			avs_readdatavalid   : out std_logic;                                        -- readdatavalid
			clock               : in  std_logic                     := 'X';             -- clk
			mem_req_address     : out std_logic_vector(25 downto 0);                    -- mem_req_address
			mem_req_byte_en     : out std_logic_vector(3 downto 0);                     -- mem_req_byte_en
			mem_req_read_writen : out std_logic;                                        -- mem_req_read_writen
			mem_req_request     : out std_logic;                                        -- mem_req_request
			mem_req_tag         : out std_logic_vector(7 downto 0);                     -- mem_req_tag
			mem_req_wdata       : out std_logic_vector(31 downto 0);                    -- mem_req_wdata
			mem_resp_dack_tag   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_resp_dack_tag
			mem_resp_data       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- mem_resp_data
			mem_resp_rack_tag   : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- mem_resp_rack_tag
		);
	end component avalon_to_mem32_bridge;

	component avalon_to_io_bridge is
		port (
			reset             : in  std_logic                     := 'X';             -- reset
			avs_read          : in  std_logic                     := 'X';             -- read
			avs_write         : in  std_logic                     := 'X';             -- write
			avs_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			avs_writedata     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			avs_ready         : out std_logic;                                        -- waitrequest_n
			avs_readdata      : out std_logic_vector(7 downto 0);                     -- readdata
			avs_readdatavalid : out std_logic;                                        -- readdatavalid
			clock             : in  std_logic                     := 'X';             -- clk
			io_ack            : in  std_logic                     := 'X';             -- ack
			io_rdata          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rdata
			io_read           : out std_logic;                                        -- read
			io_wdata          : out std_logic_vector(7 downto 0);                     -- wdata
			io_write          : out std_logic;                                        -- write
			io_address        : out std_logic_vector(19 downto 0);                    -- address
			io_irq            : in  std_logic                     := 'X';             -- irq
			avs_irq           : out std_logic                                         -- irq
		);
	end component avalon_to_io_bridge;

	component jtag_host is
		port (
			clock             : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			avs_read          : in  std_logic                     := 'X';             -- read
			avs_write         : in  std_logic                     := 'X';             -- write
			avs_address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_ready         : out std_logic;                                        -- waitrequest_n
			avs_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_readdatavalid : out std_logic;                                        -- readdatavalid
			jtag_tck          : out std_logic;                                        -- jtag_tck
			jtag_tms          : out std_logic;                                        -- jtag_tms
			jtag_tdi          : out std_logic;                                        -- jtag_tdi
			jtag_tdo          : in  std_logic                     := 'X'              -- jtag_tdo
		);
	end component jtag_host;

	component nios_tester_jtagdebug is
		port (
			mm_write_address             : out std_logic_vector(25 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_writedata           : out std_logic_vector(7 downto 0);                      -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_sink_data                 : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- data
			st_sink_valid                : in  std_logic                      := 'X';             -- valid
			st_sink_ready                : out std_logic                                          -- ready
		);
	end component nios_tester_jtagdebug;

	component nios_tester_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_tester_nios2_gen2_0;

	component nios_tester_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios_tester_onchip_memory2_0;

	component nios_tester_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_tester_pio_0;

	component nios_tester_pio_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_tester_pio_1;

	component nios_tester_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_tester_spi_0;

	component nios_tester_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			cts_n         : in  std_logic                     := 'X';             -- export
			rts_n         : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component nios_tester_uart_0;

	component nios_tester_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                      := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			audio_in_dma_mm_write_address                  : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			audio_in_dma_mm_write_waitrequest              : out std_logic;                                         -- waitrequest
			audio_in_dma_mm_write_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			audio_in_dma_mm_write_write                    : in  std_logic                      := 'X';             -- write
			audio_in_dma_mm_write_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			audio_out_dma_mm_read_address                  : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			audio_out_dma_mm_read_waitrequest              : out std_logic;                                         -- waitrequest
			audio_out_dma_mm_read_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			audio_out_dma_mm_read_read                     : in  std_logic                      := 'X';             -- read
			audio_out_dma_mm_read_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			audio_out_dma_mm_read_readdatavalid            : out std_logic;                                         -- readdatavalid
			jtagdebug_mm_write_address                     : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			jtagdebug_mm_write_waitrequest                 : out std_logic;                                         -- waitrequest
			jtagdebug_mm_write_write                       : in  std_logic                      := 'X';             -- write
			jtagdebug_mm_write_writedata                   : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_address               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                         -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                      := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                     -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                      := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                      := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                         -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                      := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                     -- readdata
			audio_in_dma_csr_address                       : out std_logic_vector(2 downto 0);                      -- address
			audio_in_dma_csr_write                         : out std_logic;                                         -- write
			audio_in_dma_csr_read                          : out std_logic;                                         -- read
			audio_in_dma_csr_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			audio_in_dma_csr_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			audio_in_dma_csr_byteenable                    : out std_logic_vector(3 downto 0);                      -- byteenable
			audio_in_dma_descriptor_slave_write            : out std_logic;                                         -- write
			audio_in_dma_descriptor_slave_writedata        : out std_logic_vector(127 downto 0);                    -- writedata
			audio_in_dma_descriptor_slave_byteenable       : out std_logic_vector(15 downto 0);                     -- byteenable
			audio_in_dma_descriptor_slave_waitrequest      : in  std_logic                      := 'X';             -- waitrequest
			audio_out_dma_csr_address                      : out std_logic_vector(2 downto 0);                      -- address
			audio_out_dma_csr_write                        : out std_logic;                                         -- write
			audio_out_dma_csr_read                         : out std_logic;                                         -- read
			audio_out_dma_csr_readdata                     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			audio_out_dma_csr_writedata                    : out std_logic_vector(31 downto 0);                     -- writedata
			audio_out_dma_csr_byteenable                   : out std_logic_vector(3 downto 0);                      -- byteenable
			audio_out_dma_descriptor_slave_write           : out std_logic;                                         -- write
			audio_out_dma_descriptor_slave_writedata       : out std_logic_vector(127 downto 0);                    -- writedata
			audio_out_dma_descriptor_slave_byteenable      : out std_logic_vector(15 downto 0);                     -- byteenable
			audio_out_dma_descriptor_slave_waitrequest     : in  std_logic                      := 'X';             -- waitrequest
			avalon2mem_0_avalon_slave_0_address            : out std_logic_vector(25 downto 0);                     -- address
			avalon2mem_0_avalon_slave_0_write              : out std_logic;                                         -- write
			avalon2mem_0_avalon_slave_0_read               : out std_logic;                                         -- read
			avalon2mem_0_avalon_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			avalon2mem_0_avalon_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			avalon2mem_0_avalon_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			avalon2mem_0_avalon_slave_0_readdatavalid      : in  std_logic                      := 'X';             -- readdatavalid
			avalon2mem_0_avalon_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			io_bridge_0_avalon_slave_0_address             : out std_logic_vector(19 downto 0);                     -- address
			io_bridge_0_avalon_slave_0_write               : out std_logic;                                         -- write
			io_bridge_0_avalon_slave_0_read                : out std_logic;                                         -- read
			io_bridge_0_avalon_slave_0_readdata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata
			io_bridge_0_avalon_slave_0_writedata           : out std_logic_vector(7 downto 0);                      -- writedata
			io_bridge_0_avalon_slave_0_readdatavalid       : in  std_logic                      := 'X';             -- readdatavalid
			io_bridge_0_avalon_slave_0_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			io_bridge_1_avalon_slave_0_address             : out std_logic_vector(19 downto 0);                     -- address
			io_bridge_1_avalon_slave_0_write               : out std_logic;                                         -- write
			io_bridge_1_avalon_slave_0_read                : out std_logic;                                         -- read
			io_bridge_1_avalon_slave_0_readdata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata
			io_bridge_1_avalon_slave_0_writedata           : out std_logic_vector(7 downto 0);                      -- writedata
			io_bridge_1_avalon_slave_0_readdatavalid       : in  std_logic                      := 'X';             -- readdatavalid
			io_bridge_1_avalon_slave_0_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			jtag_0_avalon_slave_0_address                  : out std_logic_vector(7 downto 0);                      -- address
			jtag_0_avalon_slave_0_write                    : out std_logic;                                         -- write
			jtag_0_avalon_slave_0_read                     : out std_logic;                                         -- read
			jtag_0_avalon_slave_0_readdata                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_0_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_0_avalon_slave_0_readdatavalid            : in  std_logic                      := 'X';             -- readdatavalid
			jtag_0_avalon_slave_0_waitrequest              : in  std_logic                      := 'X';             -- waitrequest
			jtag_1_avalon_slave_0_address                  : out std_logic_vector(7 downto 0);                      -- address
			jtag_1_avalon_slave_0_write                    : out std_logic;                                         -- write
			jtag_1_avalon_slave_0_read                     : out std_logic;                                         -- read
			jtag_1_avalon_slave_0_readdata                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_1_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_1_avalon_slave_0_readdatavalid            : in  std_logic                      := 'X';             -- readdatavalid
			jtag_1_avalon_slave_0_waitrequest              : in  std_logic                      := 'X';             -- waitrequest
			jtagdebug_csr_address                          : out std_logic_vector(2 downto 0);                      -- address
			jtagdebug_csr_write                            : out std_logic;                                         -- write
			jtagdebug_csr_read                             : out std_logic;                                         -- read
			jtagdebug_csr_readdata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtagdebug_csr_writedata                        : out std_logic_vector(31 downto 0);                     -- writedata
			jtagdebug_csr_byteenable                       : out std_logic_vector(3 downto 0);                      -- byteenable
			jtagdebug_descriptor_slave_write               : out std_logic;                                         -- write
			jtagdebug_descriptor_slave_writedata           : out std_logic_vector(127 downto 0);                    -- writedata
			jtagdebug_descriptor_slave_byteenable          : out std_logic_vector(15 downto 0);                     -- byteenable
			jtagdebug_descriptor_slave_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                      -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                         -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                         -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                     -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                      -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                      := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                         -- debugaccess
			onchip_memory2_0_s1_address                    : out std_logic_vector(8 downto 0);                      -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                         -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(31 downto 0);                     -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(3 downto 0);                      -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                         -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                         -- clken
			pio_0_s1_address                               : out std_logic_vector(1 downto 0);                      -- address
			pio_0_s1_write                                 : out std_logic;                                         -- write
			pio_0_s1_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			pio_0_s1_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			pio_0_s1_chipselect                            : out std_logic;                                         -- chipselect
			pio_1_s1_address                               : out std_logic_vector(2 downto 0);                      -- address
			pio_1_s1_write                                 : out std_logic;                                         -- write
			pio_1_s1_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			pio_1_s1_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			pio_1_s1_chipselect                            : out std_logic;                                         -- chipselect
			spi_0_spi_control_port_address                 : out std_logic_vector(2 downto 0);                      -- address
			spi_0_spi_control_port_write                   : out std_logic;                                         -- write
			spi_0_spi_control_port_read                    : out std_logic;                                         -- read
			spi_0_spi_control_port_readdata                : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			spi_0_spi_control_port_writedata               : out std_logic_vector(15 downto 0);                     -- writedata
			spi_0_spi_control_port_chipselect              : out std_logic;                                         -- chipselect
			uart_0_s1_address                              : out std_logic_vector(2 downto 0);                      -- address
			uart_0_s1_write                                : out std_logic;                                         -- write
			uart_0_s1_read                                 : out std_logic;                                         -- read
			uart_0_s1_readdata                             : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			uart_0_s1_writedata                            : out std_logic_vector(15 downto 0);                     -- writedata
			uart_0_s1_begintransfer                        : out std_logic;                                         -- begintransfer
			uart_0_s1_chipselect                           : out std_logic                                          -- chipselect
		);
	end component nios_tester_mm_interconnect_0;

	component nios_tester_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_tester_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_data_master_readdata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                         : std_logic;                      -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                         : std_logic;                      -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                             : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                          : std_logic_vector(3 downto 0);   -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                : std_logic;                      -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                               : std_logic;                      -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                           : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                     : std_logic_vector(31 downto 0);  -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                  : std_logic;                      -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                      : std_logic_vector(29 downto 0);  -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                         : std_logic;                      -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal audio_out_dma_mm_read_readdata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:audio_out_dma_mm_read_readdata -> audio_out_dma:mm_read_readdata
	signal audio_out_dma_mm_read_waitrequest                            : std_logic;                      -- mm_interconnect_0:audio_out_dma_mm_read_waitrequest -> audio_out_dma:mm_read_waitrequest
	signal audio_out_dma_mm_read_address                                : std_logic_vector(25 downto 0);  -- audio_out_dma:mm_read_address -> mm_interconnect_0:audio_out_dma_mm_read_address
	signal audio_out_dma_mm_read_read                                   : std_logic;                      -- audio_out_dma:mm_read_read -> mm_interconnect_0:audio_out_dma_mm_read_read
	signal audio_out_dma_mm_read_byteenable                             : std_logic_vector(3 downto 0);   -- audio_out_dma:mm_read_byteenable -> mm_interconnect_0:audio_out_dma_mm_read_byteenable
	signal audio_out_dma_mm_read_readdatavalid                          : std_logic;                      -- mm_interconnect_0:audio_out_dma_mm_read_readdatavalid -> audio_out_dma:mm_read_readdatavalid
	signal audio_in_dma_mm_write_waitrequest                            : std_logic;                      -- mm_interconnect_0:audio_in_dma_mm_write_waitrequest -> audio_in_dma:mm_write_waitrequest
	signal audio_in_dma_mm_write_address                                : std_logic_vector(25 downto 0);  -- audio_in_dma:mm_write_address -> mm_interconnect_0:audio_in_dma_mm_write_address
	signal audio_in_dma_mm_write_byteenable                             : std_logic_vector(3 downto 0);   -- audio_in_dma:mm_write_byteenable -> mm_interconnect_0:audio_in_dma_mm_write_byteenable
	signal audio_in_dma_mm_write_write                                  : std_logic;                      -- audio_in_dma:mm_write_write -> mm_interconnect_0:audio_in_dma_mm_write_write
	signal audio_in_dma_mm_write_writedata                              : std_logic_vector(31 downto 0);  -- audio_in_dma:mm_write_writedata -> mm_interconnect_0:audio_in_dma_mm_write_writedata
	signal jtagdebug_mm_write_waitrequest                               : std_logic;                      -- mm_interconnect_0:jtagdebug_mm_write_waitrequest -> jtagdebug:mm_write_waitrequest
	signal jtagdebug_mm_write_address                                   : std_logic_vector(25 downto 0);  -- jtagdebug:mm_write_address -> mm_interconnect_0:jtagdebug_mm_write_address
	signal jtagdebug_mm_write_write                                     : std_logic;                      -- jtagdebug:mm_write_write -> mm_interconnect_0:jtagdebug_mm_write_write
	signal jtagdebug_mm_write_writedata                                 : std_logic_vector(7 downto 0);   -- jtagdebug:mm_write_writedata -> mm_interconnect_0:jtagdebug_mm_write_writedata
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata        : std_logic_vector(7 downto 0);   -- io_bridge_1:avs_readdata -> mm_interconnect_0:io_bridge_1_avalon_slave_0_readdata
	signal io_bridge_1_avalon_slave_0_waitrequest                       : std_logic;                      -- io_bridge_1:avs_ready -> io_bridge_1_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_address         : std_logic_vector(19 downto 0);  -- mm_interconnect_0:io_bridge_1_avalon_slave_0_address -> io_bridge_1:avs_address
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_read            : std_logic;                      -- mm_interconnect_0:io_bridge_1_avalon_slave_0_read -> io_bridge_1:avs_read
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid   : std_logic;                      -- io_bridge_1:avs_readdatavalid -> mm_interconnect_0:io_bridge_1_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_write           : std_logic;                      -- mm_interconnect_0:io_bridge_1_avalon_slave_0_write -> io_bridge_1:avs_write
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata       : std_logic_vector(7 downto 0);   -- mm_interconnect_0:io_bridge_1_avalon_slave_0_writedata -> io_bridge_1:avs_writedata
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata       : std_logic_vector(31 downto 0);  -- avalon2mem_0:avs_readdata -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_readdata
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest    : std_logic;                      -- avalon2mem_0:avs_waitrequest -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_address        : std_logic_vector(25 downto 0);  -- mm_interconnect_0:avalon2mem_0_avalon_slave_0_address -> avalon2mem_0:avs_address
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_read           : std_logic;                      -- mm_interconnect_0:avalon2mem_0_avalon_slave_0_read -> avalon2mem_0:avs_read
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:avalon2mem_0_avalon_slave_0_byteenable -> avalon2mem_0:avs_byteenable
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid  : std_logic;                      -- avalon2mem_0:avs_readdatavalid -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_write          : std_logic;                      -- mm_interconnect_0:avalon2mem_0_avalon_slave_0_write -> avalon2mem_0:avs_write
	signal mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata      : std_logic_vector(31 downto 0);  -- mm_interconnect_0:avalon2mem_0_avalon_slave_0_writedata -> avalon2mem_0:avs_writedata
	signal mm_interconnect_0_jtag_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0);  -- jtag_0:avs_readdata -> mm_interconnect_0:jtag_0_avalon_slave_0_readdata
	signal jtag_0_avalon_slave_0_waitrequest                            : std_logic;                      -- jtag_0:avs_ready -> jtag_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_jtag_0_avalon_slave_0_address              : std_logic_vector(7 downto 0);   -- mm_interconnect_0:jtag_0_avalon_slave_0_address -> jtag_0:avs_address
	signal mm_interconnect_0_jtag_0_avalon_slave_0_read                 : std_logic;                      -- mm_interconnect_0:jtag_0_avalon_slave_0_read -> jtag_0:avs_read
	signal mm_interconnect_0_jtag_0_avalon_slave_0_readdatavalid        : std_logic;                      -- jtag_0:avs_readdatavalid -> mm_interconnect_0:jtag_0_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_jtag_0_avalon_slave_0_write                : std_logic;                      -- mm_interconnect_0:jtag_0_avalon_slave_0_write -> jtag_0:avs_write
	signal mm_interconnect_0_jtag_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_0_avalon_slave_0_writedata -> jtag_0:avs_writedata
	signal mm_interconnect_0_jtag_1_avalon_slave_0_readdata             : std_logic_vector(31 downto 0);  -- jtag_1:avs_readdata -> mm_interconnect_0:jtag_1_avalon_slave_0_readdata
	signal jtag_1_avalon_slave_0_waitrequest                            : std_logic;                      -- jtag_1:avs_ready -> jtag_1_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_jtag_1_avalon_slave_0_address              : std_logic_vector(7 downto 0);   -- mm_interconnect_0:jtag_1_avalon_slave_0_address -> jtag_1:avs_address
	signal mm_interconnect_0_jtag_1_avalon_slave_0_read                 : std_logic;                      -- mm_interconnect_0:jtag_1_avalon_slave_0_read -> jtag_1:avs_read
	signal mm_interconnect_0_jtag_1_avalon_slave_0_readdatavalid        : std_logic;                      -- jtag_1:avs_readdatavalid -> mm_interconnect_0:jtag_1_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_jtag_1_avalon_slave_0_write                : std_logic;                      -- mm_interconnect_0:jtag_1_avalon_slave_0_write -> jtag_1:avs_write
	signal mm_interconnect_0_jtag_1_avalon_slave_0_writedata            : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_1_avalon_slave_0_writedata -> jtag_1:avs_writedata
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata        : std_logic_vector(7 downto 0);   -- io_bridge_0:avs_readdata -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdata
	signal io_bridge_0_avalon_slave_0_waitrequest                       : std_logic;                      -- io_bridge_0:avs_ready -> io_bridge_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_address         : std_logic_vector(19 downto 0);  -- mm_interconnect_0:io_bridge_0_avalon_slave_0_address -> io_bridge_0:avs_address
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_read            : std_logic;                      -- mm_interconnect_0:io_bridge_0_avalon_slave_0_read -> io_bridge_0:avs_read
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid   : std_logic;                      -- io_bridge_0:avs_readdatavalid -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_write           : std_logic;                      -- mm_interconnect_0:io_bridge_0_avalon_slave_0_write -> io_bridge_0:avs_write
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata       : std_logic_vector(7 downto 0);   -- mm_interconnect_0:io_bridge_0_avalon_slave_0_writedata -> io_bridge_0:avs_writedata
	signal mm_interconnect_0_audio_out_dma_csr_readdata                 : std_logic_vector(31 downto 0);  -- audio_out_dma:csr_readdata -> mm_interconnect_0:audio_out_dma_csr_readdata
	signal mm_interconnect_0_audio_out_dma_csr_address                  : std_logic_vector(2 downto 0);   -- mm_interconnect_0:audio_out_dma_csr_address -> audio_out_dma:csr_address
	signal mm_interconnect_0_audio_out_dma_csr_read                     : std_logic;                      -- mm_interconnect_0:audio_out_dma_csr_read -> audio_out_dma:csr_read
	signal mm_interconnect_0_audio_out_dma_csr_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_0:audio_out_dma_csr_byteenable -> audio_out_dma:csr_byteenable
	signal mm_interconnect_0_audio_out_dma_csr_write                    : std_logic;                      -- mm_interconnect_0:audio_out_dma_csr_write -> audio_out_dma:csr_write
	signal mm_interconnect_0_audio_out_dma_csr_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_0:audio_out_dma_csr_writedata -> audio_out_dma:csr_writedata
	signal mm_interconnect_0_audio_in_dma_csr_readdata                  : std_logic_vector(31 downto 0);  -- audio_in_dma:csr_readdata -> mm_interconnect_0:audio_in_dma_csr_readdata
	signal mm_interconnect_0_audio_in_dma_csr_address                   : std_logic_vector(2 downto 0);   -- mm_interconnect_0:audio_in_dma_csr_address -> audio_in_dma:csr_address
	signal mm_interconnect_0_audio_in_dma_csr_read                      : std_logic;                      -- mm_interconnect_0:audio_in_dma_csr_read -> audio_in_dma:csr_read
	signal mm_interconnect_0_audio_in_dma_csr_byteenable                : std_logic_vector(3 downto 0);   -- mm_interconnect_0:audio_in_dma_csr_byteenable -> audio_in_dma:csr_byteenable
	signal mm_interconnect_0_audio_in_dma_csr_write                     : std_logic;                      -- mm_interconnect_0:audio_in_dma_csr_write -> audio_in_dma:csr_write
	signal mm_interconnect_0_audio_in_dma_csr_writedata                 : std_logic_vector(31 downto 0);  -- mm_interconnect_0:audio_in_dma_csr_writedata -> audio_in_dma:csr_writedata
	signal mm_interconnect_0_jtagdebug_csr_readdata                     : std_logic_vector(31 downto 0);  -- jtagdebug:csr_readdata -> mm_interconnect_0:jtagdebug_csr_readdata
	signal mm_interconnect_0_jtagdebug_csr_address                      : std_logic_vector(2 downto 0);   -- mm_interconnect_0:jtagdebug_csr_address -> jtagdebug:csr_address
	signal mm_interconnect_0_jtagdebug_csr_read                         : std_logic;                      -- mm_interconnect_0:jtagdebug_csr_read -> jtagdebug:csr_read
	signal mm_interconnect_0_jtagdebug_csr_byteenable                   : std_logic_vector(3 downto 0);   -- mm_interconnect_0:jtagdebug_csr_byteenable -> jtagdebug:csr_byteenable
	signal mm_interconnect_0_jtagdebug_csr_write                        : std_logic;                      -- mm_interconnect_0:jtagdebug_csr_write -> jtagdebug:csr_write
	signal mm_interconnect_0_jtagdebug_csr_writedata                    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtagdebug_csr_writedata -> jtagdebug:csr_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata      : std_logic_vector(31 downto 0);  -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest   : std_logic;                      -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess   : std_logic;                      -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address       : std_logic_vector(8 downto 0);   -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read          : std_logic;                      -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable    : std_logic_vector(3 downto 0);   -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write         : std_logic;                      -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata     : std_logic_vector(31 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_audio_out_dma_descriptor_slave_waitrequest : std_logic;                      -- audio_out_dma:descriptor_slave_waitrequest -> mm_interconnect_0:audio_out_dma_descriptor_slave_waitrequest
	signal mm_interconnect_0_audio_out_dma_descriptor_slave_byteenable  : std_logic_vector(15 downto 0);  -- mm_interconnect_0:audio_out_dma_descriptor_slave_byteenable -> audio_out_dma:descriptor_slave_byteenable
	signal mm_interconnect_0_audio_out_dma_descriptor_slave_write       : std_logic;                      -- mm_interconnect_0:audio_out_dma_descriptor_slave_write -> audio_out_dma:descriptor_slave_write
	signal mm_interconnect_0_audio_out_dma_descriptor_slave_writedata   : std_logic_vector(127 downto 0); -- mm_interconnect_0:audio_out_dma_descriptor_slave_writedata -> audio_out_dma:descriptor_slave_writedata
	signal mm_interconnect_0_audio_in_dma_descriptor_slave_waitrequest  : std_logic;                      -- audio_in_dma:descriptor_slave_waitrequest -> mm_interconnect_0:audio_in_dma_descriptor_slave_waitrequest
	signal mm_interconnect_0_audio_in_dma_descriptor_slave_byteenable   : std_logic_vector(15 downto 0);  -- mm_interconnect_0:audio_in_dma_descriptor_slave_byteenable -> audio_in_dma:descriptor_slave_byteenable
	signal mm_interconnect_0_audio_in_dma_descriptor_slave_write        : std_logic;                      -- mm_interconnect_0:audio_in_dma_descriptor_slave_write -> audio_in_dma:descriptor_slave_write
	signal mm_interconnect_0_audio_in_dma_descriptor_slave_writedata    : std_logic_vector(127 downto 0); -- mm_interconnect_0:audio_in_dma_descriptor_slave_writedata -> audio_in_dma:descriptor_slave_writedata
	signal mm_interconnect_0_jtagdebug_descriptor_slave_waitrequest     : std_logic;                      -- jtagdebug:descriptor_slave_waitrequest -> mm_interconnect_0:jtagdebug_descriptor_slave_waitrequest
	signal mm_interconnect_0_jtagdebug_descriptor_slave_byteenable      : std_logic_vector(15 downto 0);  -- mm_interconnect_0:jtagdebug_descriptor_slave_byteenable -> jtagdebug:descriptor_slave_byteenable
	signal mm_interconnect_0_jtagdebug_descriptor_slave_write           : std_logic;                      -- mm_interconnect_0:jtagdebug_descriptor_slave_write -> jtagdebug:descriptor_slave_write
	signal mm_interconnect_0_jtagdebug_descriptor_slave_writedata       : std_logic_vector(127 downto 0); -- mm_interconnect_0:jtagdebug_descriptor_slave_writedata -> jtagdebug:descriptor_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect             : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata               : std_logic_vector(31 downto 0);  -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                : std_logic_vector(8 downto 0);   -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable             : std_logic_vector(3 downto 0);   -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                  : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata              : std_logic_vector(31 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                  : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_pio_0_s1_chipselect                        : std_logic;                      -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                          : std_logic_vector(31 downto 0);  -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                             : std_logic;                      -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_0_uart_0_s1_chipselect                       : std_logic;                      -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                         : std_logic_vector(15 downto 0);  -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                             : std_logic;                      -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                    : std_logic;                      -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                            : std_logic;                      -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                        : std_logic_vector(15 downto 0);  -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal mm_interconnect_0_pio_1_s1_chipselect                        : std_logic;                      -- mm_interconnect_0:pio_1_s1_chipselect -> pio_1:chipselect
	signal mm_interconnect_0_pio_1_s1_readdata                          : std_logic_vector(31 downto 0);  -- pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	signal mm_interconnect_0_pio_1_s1_address                           : std_logic_vector(2 downto 0);   -- mm_interconnect_0:pio_1_s1_address -> pio_1:address
	signal mm_interconnect_0_pio_1_s1_write                             : std_logic;                      -- mm_interconnect_0:pio_1_s1_write -> mm_interconnect_0_pio_1_s1_write:in
	signal mm_interconnect_0_pio_1_s1_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_0:pio_1_s1_writedata -> pio_1:writedata
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect          : std_logic;                      -- mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata            : std_logic_vector(15 downto 0);  -- spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address             : std_logic_vector(2 downto 0);   -- mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                : std_logic;                      -- mm_interconnect_0:spi_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write               : std_logic;                      -- mm_interconnect_0:spi_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata           : std_logic_vector(15 downto 0);  -- mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	signal irq_mapper_receiver0_irq                                     : std_logic;                      -- audio_out_dma:csr_irq_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                     : std_logic;                      -- audio_in_dma:csr_irq_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                     : std_logic;                      -- jtagdebug:csr_irq_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                     : std_logic;                      -- io_bridge_1:avs_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                     : std_logic;                      -- pio_0:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                     : std_logic;                      -- uart_0:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                     : std_logic;                      -- spi_0:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                     : std_logic;                      -- io_bridge_0:avs_irq -> irq_mapper:receiver7_irq
	signal nios2_gen2_0_irq_irq                                         : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                               : std_logic;                      -- rst_controller:reset_out -> [avalon2mem_0:reset, io_bridge_0:reset, io_bridge_1:reset, irq_mapper:reset, jtag_0:reset, jtag_1:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                           : std_logic;                      -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal sys_reset_reset_n_ports_inv                                  : std_logic;                      -- sys_reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_io_bridge_1_avalon_slave_0_inv             : std_logic;                      -- io_bridge_1_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:io_bridge_1_avalon_slave_0_waitrequest
	signal mm_interconnect_0_jtag_0_avalon_slave_0_inv                  : std_logic;                      -- jtag_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:jtag_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_jtag_1_avalon_slave_0_inv                  : std_logic;                      -- jtag_1_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:jtag_1_avalon_slave_0_waitrequest
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_inv             : std_logic;                      -- io_bridge_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:io_bridge_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                   : std_logic;                      -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv                   : std_logic;                      -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv                  : std_logic;                      -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal mm_interconnect_0_pio_1_s1_write_ports_inv                   : std_logic;                      -- mm_interconnect_0_pio_1_s1_write:inv -> pio_1:write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv      : std_logic;                      -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> spi_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv     : std_logic;                      -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> spi_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                      -- rst_controller_reset_out_reset:inv -> [audio_in_dma:reset_n_reset_n, audio_out_dma:reset_n_reset_n, jtagdebug:reset_n_reset_n, nios2_gen2_0:reset_n, pio_0:reset_n, pio_1:reset_n, spi_0:reset_n, uart_0:reset_n]

begin

	audio_in_dma : component nios_tester_audio_in_dma
		port map (
			mm_write_address             => audio_in_dma_mm_write_address,                               --         mm_write.address
			mm_write_write               => audio_in_dma_mm_write_write,                                 --                 .write
			mm_write_byteenable          => audio_in_dma_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => audio_in_dma_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => audio_in_dma_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => sys_clock_clk,                                               --            clock.clk
			reset_n_reset_n              => rst_controller_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_audio_in_dma_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_audio_in_dma_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_audio_in_dma_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_audio_in_dma_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_audio_in_dma_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_audio_in_dma_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_audio_in_dma_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_audio_in_dma_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_audio_in_dma_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_audio_in_dma_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver1_irq,                                    --          csr_irq.irq
			st_sink_data                 => audio_in_data,                                               --          st_sink.data
			st_sink_valid                => audio_in_valid,                                              --                 .valid
			st_sink_ready                => audio_in_ready                                               --                 .ready
		);

	audio_out_dma : component nios_tester_audio_out_dma
		port map (
			mm_read_address              => audio_out_dma_mm_read_address,                                --          mm_read.address
			mm_read_read                 => audio_out_dma_mm_read_read,                                   --                 .read
			mm_read_byteenable           => audio_out_dma_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => audio_out_dma_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => audio_out_dma_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => audio_out_dma_mm_read_readdatavalid,                          --                 .readdatavalid
			clock_clk                    => sys_clock_clk,                                                --            clock.clk
			reset_n_reset_n              => rst_controller_reset_out_reset_ports_inv,                     --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_audio_out_dma_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_audio_out_dma_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_audio_out_dma_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_audio_out_dma_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_audio_out_dma_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_audio_out_dma_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_audio_out_dma_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_audio_out_dma_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_audio_out_dma_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_audio_out_dma_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver0_irq,                                     --          csr_irq.irq
			st_source_data               => audio_out_data,                                               --        st_source.data
			st_source_valid              => audio_out_valid,                                              --                 .valid
			st_source_ready              => audio_out_ready                                               --                 .ready
		);

	avalon2mem_0 : component avalon_to_mem32_bridge
		generic map (
			g_tag => "01011011"
		)
		port map (
			reset               => rst_controller_reset_out_reset,                              --          reset.reset
			avs_read            => mm_interconnect_0_avalon2mem_0_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write           => mm_interconnect_0_avalon2mem_0_avalon_slave_0_write,         --               .write
			avs_address         => mm_interconnect_0_avalon2mem_0_avalon_slave_0_address,       --               .address
			avs_writedata       => mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata,     --               .writedata
			avs_byteenable      => mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable,    --               .byteenable
			avs_waitrequest     => mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest,   --               .waitrequest
			avs_readdata        => mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid   => mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid, --               .readdatavalid
			clock               => sys_clock_clk,                                               --          clock.clk
			mem_req_address     => mem_mem_req_address,                                         --            mem.mem_req_address
			mem_req_byte_en     => mem_mem_req_byte_en,                                         --               .mem_req_byte_en
			mem_req_read_writen => mem_mem_req_read_writen,                                     --               .mem_req_read_writen
			mem_req_request     => mem_mem_req_request,                                         --               .mem_req_request
			mem_req_tag         => mem_mem_req_tag,                                             --               .mem_req_tag
			mem_req_wdata       => mem_mem_req_wdata,                                           --               .mem_req_wdata
			mem_resp_dack_tag   => mem_mem_resp_dack_tag,                                       --               .mem_resp_dack_tag
			mem_resp_data       => mem_mem_resp_data,                                           --               .mem_resp_data
			mem_resp_rack_tag   => mem_mem_resp_rack_tag                                        --               .mem_resp_rack_tag
		);

	io_bridge_0 : component avalon_to_io_bridge
		port map (
			reset             => rst_controller_reset_out_reset,                             --          reset.reset
			avs_read          => mm_interconnect_0_io_bridge_0_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write         => mm_interconnect_0_io_bridge_0_avalon_slave_0_write,         --               .write
			avs_address       => mm_interconnect_0_io_bridge_0_avalon_slave_0_address,       --               .address
			avs_writedata     => mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata,     --               .writedata
			avs_ready         => io_bridge_0_avalon_slave_0_waitrequest,                     --               .waitrequest_n
			avs_readdata      => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid, --               .readdatavalid
			clock             => sys_clock_clk,                                              --          clock.clk
			io_ack            => io_ack,                                                     --             io.ack
			io_rdata          => io_rdata,                                                   --               .rdata
			io_read           => io_read,                                                    --               .read
			io_wdata          => io_wdata,                                                   --               .wdata
			io_write          => io_write,                                                   --               .write
			io_address        => io_address,                                                 --               .address
			io_irq            => io_irq,                                                     --               .irq
			avs_irq           => irq_mapper_receiver7_irq                                    --            irq.irq
		);

	io_bridge_1 : component avalon_to_io_bridge
		port map (
			reset             => rst_controller_reset_out_reset,                             --          reset.reset
			avs_read          => mm_interconnect_0_io_bridge_1_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write         => mm_interconnect_0_io_bridge_1_avalon_slave_0_write,         --               .write
			avs_address       => mm_interconnect_0_io_bridge_1_avalon_slave_0_address,       --               .address
			avs_writedata     => mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata,     --               .writedata
			avs_ready         => io_bridge_1_avalon_slave_0_waitrequest,                     --               .waitrequest_n
			avs_readdata      => mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid => mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid, --               .readdatavalid
			clock             => sys_clock_clk,                                              --          clock.clk
			io_ack            => io_u2p_ack,                                                 --             io.ack
			io_rdata          => io_u2p_rdata,                                               --               .rdata
			io_read           => io_u2p_read,                                                --               .read
			io_wdata          => io_u2p_wdata,                                               --               .wdata
			io_write          => io_u2p_write,                                               --               .write
			io_address        => io_u2p_address,                                             --               .address
			io_irq            => io_u2p_irq,                                                 --               .irq
			avs_irq           => irq_mapper_receiver3_irq                                    --            irq.irq
		);

	jtag_0 : component jtag_host
		port map (
			clock             => sys_clock_clk,                                         --          clock.clk
			reset             => rst_controller_reset_out_reset,                        --          reset.reset
			avs_read          => mm_interconnect_0_jtag_0_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write         => mm_interconnect_0_jtag_0_avalon_slave_0_write,         --               .write
			avs_address       => mm_interconnect_0_jtag_0_avalon_slave_0_address,       --               .address
			avs_writedata     => mm_interconnect_0_jtag_0_avalon_slave_0_writedata,     --               .writedata
			avs_ready         => jtag_0_avalon_slave_0_waitrequest,                     --               .waitrequest_n
			avs_readdata      => mm_interconnect_0_jtag_0_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid => mm_interconnect_0_jtag_0_avalon_slave_0_readdatavalid, --               .readdatavalid
			jtag_tck          => jtag0_jtag_tck,                                        --           jtag.jtag_tck
			jtag_tms          => jtag0_jtag_tms,                                        --               .jtag_tms
			jtag_tdi          => jtag0_jtag_tdi,                                        --               .jtag_tdi
			jtag_tdo          => jtag0_jtag_tdo                                         --               .jtag_tdo
		);

	jtag_1 : component jtag_host
		port map (
			clock             => sys_clock_clk,                                         --          clock.clk
			reset             => rst_controller_reset_out_reset,                        --          reset.reset
			avs_read          => mm_interconnect_0_jtag_1_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write         => mm_interconnect_0_jtag_1_avalon_slave_0_write,         --               .write
			avs_address       => mm_interconnect_0_jtag_1_avalon_slave_0_address,       --               .address
			avs_writedata     => mm_interconnect_0_jtag_1_avalon_slave_0_writedata,     --               .writedata
			avs_ready         => jtag_1_avalon_slave_0_waitrequest,                     --               .waitrequest_n
			avs_readdata      => mm_interconnect_0_jtag_1_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid => mm_interconnect_0_jtag_1_avalon_slave_0_readdatavalid, --               .readdatavalid
			jtag_tck          => jtag1_jtag_tck,                                        --           jtag.jtag_tck
			jtag_tms          => jtag1_jtag_tms,                                        --               .jtag_tms
			jtag_tdi          => jtag1_jtag_tdi,                                        --               .jtag_tdi
			jtag_tdo          => jtag1_jtag_tdo                                         --               .jtag_tdo
		);

	jtagdebug : component nios_tester_jtagdebug
		port map (
			mm_write_address             => jtagdebug_mm_write_address,                               --         mm_write.address
			mm_write_write               => jtagdebug_mm_write_write,                                 --                 .write
			mm_write_writedata           => jtagdebug_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => jtagdebug_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => sys_clock_clk,                                            --            clock.clk
			reset_n_reset_n              => rst_controller_reset_out_reset_ports_inv,                 --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_jtagdebug_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_jtagdebug_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_jtagdebug_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_jtagdebug_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_jtagdebug_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_jtagdebug_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_jtagdebug_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_jtagdebug_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_jtagdebug_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_jtagdebug_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver2_irq,                                 --          csr_irq.irq
			st_sink_data                 => jtag_in_data,                                             --          st_sink.data
			st_sink_valid                => jtag_in_valid,                                            --                 .valid
			st_sink_ready                => jtag_in_ready                                             --                 .ready
		);

	nios2_gen2_0 : component nios_tester_nios2_gen2_0
		port map (
			clk                                 => sys_clock_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component nios_tester_onchip_memory2_0
		port map (
			clk        => sys_clock_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	pio_0 : component nios_tester_pio_0
		port map (
			clk        => sys_clock_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			in_port    => dummy_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                    --                 irq.irq
		);

	pio_1 : component nios_tester_pio_1
		port map (
			clk        => sys_clock_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_1_s1_readdata,        --                    .readdata
			in_port    => pio_in_port,                                -- external_connection.export
			out_port   => pio_out_port                                --                    .export
		);

	spi_0 : component nios_tester_spi_0
		port map (
			clk           => sys_clock_clk,                                            --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver6_irq,                                 --              irq.irq
			MISO          => spi_MISO,                                                 --         external.export
			MOSI          => spi_MOSI,                                                 --                 .export
			SCLK          => spi_SCLK,                                                 --                 .export
			SS_n          => spi_SS_n                                                  --                 .export
		);

	uart_0 : component nios_tester_uart_0
		port map (
			clk           => sys_clock_clk,                               --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			dataavailable => open,                                        --                    .dataavailable
			readyfordata  => open,                                        --                    .readyfordata
			rxd           => uart_rxd,                                    -- external_connection.export
			txd           => uart_txd,                                    --                    .export
			cts_n         => uart_cts_n,                                  --                    .export
			rts_n         => uart_rts_n,                                  --                    .export
			irq           => irq_mapper_receiver5_irq                     --                 irq.irq
		);

	mm_interconnect_0 : component nios_tester_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => sys_clock_clk,                                                --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                               -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			audio_in_dma_mm_write_address                  => audio_in_dma_mm_write_address,                                --                    audio_in_dma_mm_write.address
			audio_in_dma_mm_write_waitrequest              => audio_in_dma_mm_write_waitrequest,                            --                                         .waitrequest
			audio_in_dma_mm_write_byteenable               => audio_in_dma_mm_write_byteenable,                             --                                         .byteenable
			audio_in_dma_mm_write_write                    => audio_in_dma_mm_write_write,                                  --                                         .write
			audio_in_dma_mm_write_writedata                => audio_in_dma_mm_write_writedata,                              --                                         .writedata
			audio_out_dma_mm_read_address                  => audio_out_dma_mm_read_address,                                --                    audio_out_dma_mm_read.address
			audio_out_dma_mm_read_waitrequest              => audio_out_dma_mm_read_waitrequest,                            --                                         .waitrequest
			audio_out_dma_mm_read_byteenable               => audio_out_dma_mm_read_byteenable,                             --                                         .byteenable
			audio_out_dma_mm_read_read                     => audio_out_dma_mm_read_read,                                   --                                         .read
			audio_out_dma_mm_read_readdata                 => audio_out_dma_mm_read_readdata,                               --                                         .readdata
			audio_out_dma_mm_read_readdatavalid            => audio_out_dma_mm_read_readdatavalid,                          --                                         .readdatavalid
			jtagdebug_mm_write_address                     => jtagdebug_mm_write_address,                                   --                       jtagdebug_mm_write.address
			jtagdebug_mm_write_waitrequest                 => jtagdebug_mm_write_waitrequest,                               --                                         .waitrequest
			jtagdebug_mm_write_write                       => jtagdebug_mm_write_write,                                     --                                         .write
			jtagdebug_mm_write_writedata                   => jtagdebug_mm_write_writedata,                                 --                                         .writedata
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                             --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                         --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                          --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                                --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                            --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                               --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                           --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                         --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                      --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                  --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                         --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                     --                                         .readdata
			audio_in_dma_csr_address                       => mm_interconnect_0_audio_in_dma_csr_address,                   --                         audio_in_dma_csr.address
			audio_in_dma_csr_write                         => mm_interconnect_0_audio_in_dma_csr_write,                     --                                         .write
			audio_in_dma_csr_read                          => mm_interconnect_0_audio_in_dma_csr_read,                      --                                         .read
			audio_in_dma_csr_readdata                      => mm_interconnect_0_audio_in_dma_csr_readdata,                  --                                         .readdata
			audio_in_dma_csr_writedata                     => mm_interconnect_0_audio_in_dma_csr_writedata,                 --                                         .writedata
			audio_in_dma_csr_byteenable                    => mm_interconnect_0_audio_in_dma_csr_byteenable,                --                                         .byteenable
			audio_in_dma_descriptor_slave_write            => mm_interconnect_0_audio_in_dma_descriptor_slave_write,        --            audio_in_dma_descriptor_slave.write
			audio_in_dma_descriptor_slave_writedata        => mm_interconnect_0_audio_in_dma_descriptor_slave_writedata,    --                                         .writedata
			audio_in_dma_descriptor_slave_byteenable       => mm_interconnect_0_audio_in_dma_descriptor_slave_byteenable,   --                                         .byteenable
			audio_in_dma_descriptor_slave_waitrequest      => mm_interconnect_0_audio_in_dma_descriptor_slave_waitrequest,  --                                         .waitrequest
			audio_out_dma_csr_address                      => mm_interconnect_0_audio_out_dma_csr_address,                  --                        audio_out_dma_csr.address
			audio_out_dma_csr_write                        => mm_interconnect_0_audio_out_dma_csr_write,                    --                                         .write
			audio_out_dma_csr_read                         => mm_interconnect_0_audio_out_dma_csr_read,                     --                                         .read
			audio_out_dma_csr_readdata                     => mm_interconnect_0_audio_out_dma_csr_readdata,                 --                                         .readdata
			audio_out_dma_csr_writedata                    => mm_interconnect_0_audio_out_dma_csr_writedata,                --                                         .writedata
			audio_out_dma_csr_byteenable                   => mm_interconnect_0_audio_out_dma_csr_byteenable,               --                                         .byteenable
			audio_out_dma_descriptor_slave_write           => mm_interconnect_0_audio_out_dma_descriptor_slave_write,       --           audio_out_dma_descriptor_slave.write
			audio_out_dma_descriptor_slave_writedata       => mm_interconnect_0_audio_out_dma_descriptor_slave_writedata,   --                                         .writedata
			audio_out_dma_descriptor_slave_byteenable      => mm_interconnect_0_audio_out_dma_descriptor_slave_byteenable,  --                                         .byteenable
			audio_out_dma_descriptor_slave_waitrequest     => mm_interconnect_0_audio_out_dma_descriptor_slave_waitrequest, --                                         .waitrequest
			avalon2mem_0_avalon_slave_0_address            => mm_interconnect_0_avalon2mem_0_avalon_slave_0_address,        --              avalon2mem_0_avalon_slave_0.address
			avalon2mem_0_avalon_slave_0_write              => mm_interconnect_0_avalon2mem_0_avalon_slave_0_write,          --                                         .write
			avalon2mem_0_avalon_slave_0_read               => mm_interconnect_0_avalon2mem_0_avalon_slave_0_read,           --                                         .read
			avalon2mem_0_avalon_slave_0_readdata           => mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata,       --                                         .readdata
			avalon2mem_0_avalon_slave_0_writedata          => mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata,      --                                         .writedata
			avalon2mem_0_avalon_slave_0_byteenable         => mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable,     --                                         .byteenable
			avalon2mem_0_avalon_slave_0_readdatavalid      => mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid,  --                                         .readdatavalid
			avalon2mem_0_avalon_slave_0_waitrequest        => mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest,    --                                         .waitrequest
			io_bridge_0_avalon_slave_0_address             => mm_interconnect_0_io_bridge_0_avalon_slave_0_address,         --               io_bridge_0_avalon_slave_0.address
			io_bridge_0_avalon_slave_0_write               => mm_interconnect_0_io_bridge_0_avalon_slave_0_write,           --                                         .write
			io_bridge_0_avalon_slave_0_read                => mm_interconnect_0_io_bridge_0_avalon_slave_0_read,            --                                         .read
			io_bridge_0_avalon_slave_0_readdata            => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata,        --                                         .readdata
			io_bridge_0_avalon_slave_0_writedata           => mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata,       --                                         .writedata
			io_bridge_0_avalon_slave_0_readdatavalid       => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid,   --                                         .readdatavalid
			io_bridge_0_avalon_slave_0_waitrequest         => mm_interconnect_0_io_bridge_0_avalon_slave_0_inv,             --                                         .waitrequest
			io_bridge_1_avalon_slave_0_address             => mm_interconnect_0_io_bridge_1_avalon_slave_0_address,         --               io_bridge_1_avalon_slave_0.address
			io_bridge_1_avalon_slave_0_write               => mm_interconnect_0_io_bridge_1_avalon_slave_0_write,           --                                         .write
			io_bridge_1_avalon_slave_0_read                => mm_interconnect_0_io_bridge_1_avalon_slave_0_read,            --                                         .read
			io_bridge_1_avalon_slave_0_readdata            => mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata,        --                                         .readdata
			io_bridge_1_avalon_slave_0_writedata           => mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata,       --                                         .writedata
			io_bridge_1_avalon_slave_0_readdatavalid       => mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid,   --                                         .readdatavalid
			io_bridge_1_avalon_slave_0_waitrequest         => mm_interconnect_0_io_bridge_1_avalon_slave_0_inv,             --                                         .waitrequest
			jtag_0_avalon_slave_0_address                  => mm_interconnect_0_jtag_0_avalon_slave_0_address,              --                    jtag_0_avalon_slave_0.address
			jtag_0_avalon_slave_0_write                    => mm_interconnect_0_jtag_0_avalon_slave_0_write,                --                                         .write
			jtag_0_avalon_slave_0_read                     => mm_interconnect_0_jtag_0_avalon_slave_0_read,                 --                                         .read
			jtag_0_avalon_slave_0_readdata                 => mm_interconnect_0_jtag_0_avalon_slave_0_readdata,             --                                         .readdata
			jtag_0_avalon_slave_0_writedata                => mm_interconnect_0_jtag_0_avalon_slave_0_writedata,            --                                         .writedata
			jtag_0_avalon_slave_0_readdatavalid            => mm_interconnect_0_jtag_0_avalon_slave_0_readdatavalid,        --                                         .readdatavalid
			jtag_0_avalon_slave_0_waitrequest              => mm_interconnect_0_jtag_0_avalon_slave_0_inv,                  --                                         .waitrequest
			jtag_1_avalon_slave_0_address                  => mm_interconnect_0_jtag_1_avalon_slave_0_address,              --                    jtag_1_avalon_slave_0.address
			jtag_1_avalon_slave_0_write                    => mm_interconnect_0_jtag_1_avalon_slave_0_write,                --                                         .write
			jtag_1_avalon_slave_0_read                     => mm_interconnect_0_jtag_1_avalon_slave_0_read,                 --                                         .read
			jtag_1_avalon_slave_0_readdata                 => mm_interconnect_0_jtag_1_avalon_slave_0_readdata,             --                                         .readdata
			jtag_1_avalon_slave_0_writedata                => mm_interconnect_0_jtag_1_avalon_slave_0_writedata,            --                                         .writedata
			jtag_1_avalon_slave_0_readdatavalid            => mm_interconnect_0_jtag_1_avalon_slave_0_readdatavalid,        --                                         .readdatavalid
			jtag_1_avalon_slave_0_waitrequest              => mm_interconnect_0_jtag_1_avalon_slave_0_inv,                  --                                         .waitrequest
			jtagdebug_csr_address                          => mm_interconnect_0_jtagdebug_csr_address,                      --                            jtagdebug_csr.address
			jtagdebug_csr_write                            => mm_interconnect_0_jtagdebug_csr_write,                        --                                         .write
			jtagdebug_csr_read                             => mm_interconnect_0_jtagdebug_csr_read,                         --                                         .read
			jtagdebug_csr_readdata                         => mm_interconnect_0_jtagdebug_csr_readdata,                     --                                         .readdata
			jtagdebug_csr_writedata                        => mm_interconnect_0_jtagdebug_csr_writedata,                    --                                         .writedata
			jtagdebug_csr_byteenable                       => mm_interconnect_0_jtagdebug_csr_byteenable,                   --                                         .byteenable
			jtagdebug_descriptor_slave_write               => mm_interconnect_0_jtagdebug_descriptor_slave_write,           --               jtagdebug_descriptor_slave.write
			jtagdebug_descriptor_slave_writedata           => mm_interconnect_0_jtagdebug_descriptor_slave_writedata,       --                                         .writedata
			jtagdebug_descriptor_slave_byteenable          => mm_interconnect_0_jtagdebug_descriptor_slave_byteenable,      --                                         .byteenable
			jtagdebug_descriptor_slave_waitrequest         => mm_interconnect_0_jtagdebug_descriptor_slave_waitrequest,     --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,       --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,         --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,          --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,      --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,     --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,    --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,   --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,   --                                         .debugaccess
			onchip_memory2_0_s1_address                    => mm_interconnect_0_onchip_memory2_0_s1_address,                --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_0_onchip_memory2_0_s1_write,                  --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,               --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,              --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,             --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,             --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                  --                                         .clken
			pio_0_s1_address                               => mm_interconnect_0_pio_0_s1_address,                           --                                 pio_0_s1.address
			pio_0_s1_write                                 => mm_interconnect_0_pio_0_s1_write,                             --                                         .write
			pio_0_s1_readdata                              => mm_interconnect_0_pio_0_s1_readdata,                          --                                         .readdata
			pio_0_s1_writedata                             => mm_interconnect_0_pio_0_s1_writedata,                         --                                         .writedata
			pio_0_s1_chipselect                            => mm_interconnect_0_pio_0_s1_chipselect,                        --                                         .chipselect
			pio_1_s1_address                               => mm_interconnect_0_pio_1_s1_address,                           --                                 pio_1_s1.address
			pio_1_s1_write                                 => mm_interconnect_0_pio_1_s1_write,                             --                                         .write
			pio_1_s1_readdata                              => mm_interconnect_0_pio_1_s1_readdata,                          --                                         .readdata
			pio_1_s1_writedata                             => mm_interconnect_0_pio_1_s1_writedata,                         --                                         .writedata
			pio_1_s1_chipselect                            => mm_interconnect_0_pio_1_s1_chipselect,                        --                                         .chipselect
			spi_0_spi_control_port_address                 => mm_interconnect_0_spi_0_spi_control_port_address,             --                   spi_0_spi_control_port.address
			spi_0_spi_control_port_write                   => mm_interconnect_0_spi_0_spi_control_port_write,               --                                         .write
			spi_0_spi_control_port_read                    => mm_interconnect_0_spi_0_spi_control_port_read,                --                                         .read
			spi_0_spi_control_port_readdata                => mm_interconnect_0_spi_0_spi_control_port_readdata,            --                                         .readdata
			spi_0_spi_control_port_writedata               => mm_interconnect_0_spi_0_spi_control_port_writedata,           --                                         .writedata
			spi_0_spi_control_port_chipselect              => mm_interconnect_0_spi_0_spi_control_port_chipselect,          --                                         .chipselect
			uart_0_s1_address                              => mm_interconnect_0_uart_0_s1_address,                          --                                uart_0_s1.address
			uart_0_s1_write                                => mm_interconnect_0_uart_0_s1_write,                            --                                         .write
			uart_0_s1_read                                 => mm_interconnect_0_uart_0_s1_read,                             --                                         .read
			uart_0_s1_readdata                             => mm_interconnect_0_uart_0_s1_readdata,                         --                                         .readdata
			uart_0_s1_writedata                            => mm_interconnect_0_uart_0_s1_writedata,                        --                                         .writedata
			uart_0_s1_begintransfer                        => mm_interconnect_0_uart_0_s1_begintransfer,                    --                                         .begintransfer
			uart_0_s1_chipselect                           => mm_interconnect_0_uart_0_s1_chipselect                        --                                         .chipselect
		);

	irq_mapper : component nios_tester_irq_mapper
		port map (
			clk           => sys_clock_clk,                  --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,       -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,       -- receiver7.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => sys_clock_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

	mm_interconnect_0_io_bridge_1_avalon_slave_0_inv <= not io_bridge_1_avalon_slave_0_waitrequest;

	mm_interconnect_0_jtag_0_avalon_slave_0_inv <= not jtag_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_jtag_1_avalon_slave_0_inv <= not jtag_1_avalon_slave_0_waitrequest;

	mm_interconnect_0_io_bridge_0_avalon_slave_0_inv <= not io_bridge_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	mm_interconnect_0_pio_1_s1_write_ports_inv <= not mm_interconnect_0_pio_1_s1_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_tester
