
library ieee;
use ieee.std_logic_1164.all;

entity mk7_pla is
port (
    A       : in  std_logic_vector(7 downto 0);
    Q       : out std_logic_vector(4 downto 1) );
end mk7_pla;

architecture table of mk7_pla is
begin
    process(A)
    begin
        Q <= X"F";
        if A(7)='0' then
            Q <= "101" & not A(3);
        else
            case A(6 downto 0) is
                when "0000000" => Q <= "0110";
                when "0000001" => Q <= "0111";
                when "0000010" => Q <= "1111";
                when "0000011" => Q <= "1111";
                when "0000100" => Q <= "0010";
                when "0000101" => Q <= "0011";
                when "0000110" => Q <= "1010";
                when "0000111" => Q <= "1011";
                when "0001000" => Q <= "0110";
                when "0001001" => Q <= "0111";
                when "0001010" => Q <= "1111";
                when "0001011" => Q <= "1111";
                when "0001100" => Q <= "0010";
                when "0001101" => Q <= "0011";
                when "0001110" => Q <= "1010";
                when "0001111" => Q <= "1011";
                when "0010000" => Q <= "0110";
                when "0010001" => Q <= "0111";
                when "0010010" => Q <= "1111";
                when "0010011" => Q <= "1111";
                when "0010100" => Q <= "0010";
                when "0010101" => Q <= "0011";
                when "0010110" => Q <= "1010";
                when "0010111" => Q <= "1011";
                when "0011000" => Q <= "0110";
                when "0011001" => Q <= "0111";
                when "0011010" => Q <= "1111";
                when "0011011" => Q <= "1111";
                when "0011100" => Q <= "0010";
                when "0011101" => Q <= "0011";
                when "0011110" => Q <= "1010";
                when "0011111" => Q <= "1011";
                when "0100000" => Q <= "0110";
                when "0100001" => Q <= "0111";
                when "0100010" => Q <= "1111";
                when "0100011" => Q <= "1111";
                when "0100100" => Q <= "0010";
                when "0100101" => Q <= "0011";
                when "0100110" => Q <= "1010";
                when "0100111" => Q <= "1011";
                when "0101000" => Q <= "0110";
                when "0101001" => Q <= "0101";
                when "0101010" => Q <= "1111";
                when "0101011" => Q <= "1101";
                when "0101100" => Q <= "0011";
                when "0101101" => Q <= "0001";
                when "0101110" => Q <= "1010";
                when "0101111" => Q <= "1001";
                when "0110000" => Q <= "0111";
                when "0110001" => Q <= "0111";
                when "0110010" => Q <= "1111";
                when "0110011" => Q <= "1111";
                when "0110100" => Q <= "0011";
                when "0110101" => Q <= "0011";
                when "0110110" => Q <= "1010";
                when "0110111" => Q <= "1010";
                when "0111000" => Q <= "0111";
                when "0111001" => Q <= "0111";
                when "0111010" => Q <= "1111";
                when "0111011" => Q <= "1111";
                when "0111100" => Q <= "0010";
                when "0111101" => Q <= "0010";
                when "0111110" => Q <= "1011";
                when "0111111" => Q <= "1010";
                when "1000000" => Q <= "0110";
                when "1000001" => Q <= "0111";
                when "1000010" => Q <= "1111";
                when "1000011" => Q <= "1111";
                when "1000100" => Q <= "0010";
                when "1000101" => Q <= "0011";
                when "1000110" => Q <= "1010";
                when "1000111" => Q <= "1011";
                when "1001000" => Q <= "0110";
                when "1001001" => Q <= "0111";
                when "1001010" => Q <= "1111";
                when "1001011" => Q <= "1111";
                when "1001100" => Q <= "0010";
                when "1001101" => Q <= "0011";
                when "1001110" => Q <= "1010";
                when "1001111" => Q <= "1011";
                when "1010000" => Q <= "0110";
                when "1010001" => Q <= "0111";
                when "1010010" => Q <= "1111";
                when "1010011" => Q <= "1111";
                when "1010100" => Q <= "0010";
                when "1010101" => Q <= "0011";
                when "1010110" => Q <= "1010";
                when "1010111" => Q <= "1011";
                when "1011000" => Q <= "0110";
                when "1011001" => Q <= "0111";
                when "1011010" => Q <= "1111";
                when "1011011" => Q <= "1111";
                when "1011100" => Q <= "0010";
                when "1011101" => Q <= "0011";
                when "1011110" => Q <= "1010";
                when "1011111" => Q <= "1011";
                when "1100000" => Q <= "0110";
                when "1100001" => Q <= "0101";
                when "1100010" => Q <= "1110";
                when "1100011" => Q <= "1101";
                when "1100100" => Q <= "0011";
                when "1100101" => Q <= "0001";
                when "1100110" => Q <= "1011";
                when "1100111" => Q <= "1001";
                when "1101000" => Q <= "0111";
                when "1101001" => Q <= "0111";
                when "1101010" => Q <= "1111";
                when "1101011" => Q <= "1111";
                when "1101100" => Q <= "0011";
                when "1101101" => Q <= "0011";
                when "1101110" => Q <= "1011";
                when "1101111" => Q <= "1011";
                when "1110000" => Q <= "0111";
                when "1110001" => Q <= "0111";
                when "1110010" => Q <= "1111";
                when "1110011" => Q <= "1111";
                when "1110100" => Q <= "0011";
                when "1110101" => Q <= "0011";
                when "1110110" => Q <= "1010";
                when "1110111" => Q <= "1010";
                when "1111000" => Q <= "0111";
                when "1111001" => Q <= "0111";
                when "1111010" => Q <= "1111";
                when "1111011" => Q <= "1111";
                when "1111100" => Q <= "0011";
                when "1111101" => Q <= "0011";
                when "1111110" => Q <= "1010";
                when "1111111" => Q <= "1010";
                when others    => Q <= "1111";
            end case;
        end if;            
    end process;
end table;
