// nios_solo.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module nios_solo (
		input  wire        clk_clk,                 //    clk.clk
		input  wire        io_ack,                  //     io.ack
		input  wire [7:0]  io_rdata,                //       .rdata
		output wire        io_read,                 //       .read
		output wire [7:0]  io_wdata,                //       .wdata
		output wire        io_write,                //       .write
		output wire [19:0] io_address,              //       .address
		input  wire        io_irq,                  //       .irq
		input  wire        io_u2p_ack,              // io_u2p.ack
		input  wire [7:0]  io_u2p_rdata,            //       .rdata
		output wire        io_u2p_read,             //       .read
		output wire [7:0]  io_u2p_wdata,            //       .wdata
		output wire        io_u2p_write,            //       .write
		output wire [19:0] io_u2p_address,          //       .address
		input  wire        io_u2p_irq,              //       .irq
		output wire [25:0] mem_mem_req_address,     //    mem.mem_req_address
		output wire [3:0]  mem_mem_req_byte_en,     //       .mem_req_byte_en
		output wire        mem_mem_req_read_writen, //       .mem_req_read_writen
		output wire        mem_mem_req_request,     //       .mem_req_request
		output wire [7:0]  mem_mem_req_tag,         //       .mem_req_tag
		output wire [31:0] mem_mem_req_wdata,       //       .mem_req_wdata
		input  wire [7:0]  mem_mem_resp_dack_tag,   //       .mem_resp_dack_tag
		input  wire [31:0] mem_mem_resp_data,       //       .mem_resp_data
		input  wire [7:0]  mem_mem_resp_rack_tag,   //       .mem_resp_rack_tag
		input  wire        reset_reset_n            //  reset.reset_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [31:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [29:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire   [7:0] mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata;       // io_bridge_0:avs_readdata -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_io_bridge_0_avalon_slave_0_waitrequest;    // io_bridge_0:avs_ready -> mm_interconnect_0:io_bridge_0_avalon_slave_0_waitrequest
	wire  [19:0] mm_interconnect_0_io_bridge_0_avalon_slave_0_address;        // mm_interconnect_0:io_bridge_0_avalon_slave_0_address -> io_bridge_0:avs_address
	wire         mm_interconnect_0_io_bridge_0_avalon_slave_0_read;           // mm_interconnect_0:io_bridge_0_avalon_slave_0_read -> io_bridge_0:avs_read
	wire         mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid;  // io_bridge_0:avs_readdatavalid -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_io_bridge_0_avalon_slave_0_write;          // mm_interconnect_0:io_bridge_0_avalon_slave_0_write -> io_bridge_0:avs_write
	wire   [7:0] mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata;      // mm_interconnect_0:io_bridge_0_avalon_slave_0_writedata -> io_bridge_0:avs_writedata
	wire   [7:0] mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata;       // io_bridge_1:avs_readdata -> mm_interconnect_0:io_bridge_1_avalon_slave_0_readdata
	wire         mm_interconnect_0_io_bridge_1_avalon_slave_0_waitrequest;    // io_bridge_1:avs_ready -> mm_interconnect_0:io_bridge_1_avalon_slave_0_waitrequest
	wire  [19:0] mm_interconnect_0_io_bridge_1_avalon_slave_0_address;        // mm_interconnect_0:io_bridge_1_avalon_slave_0_address -> io_bridge_1:avs_address
	wire         mm_interconnect_0_io_bridge_1_avalon_slave_0_read;           // mm_interconnect_0:io_bridge_1_avalon_slave_0_read -> io_bridge_1:avs_read
	wire         mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid;  // io_bridge_1:avs_readdatavalid -> mm_interconnect_0:io_bridge_1_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_io_bridge_1_avalon_slave_0_write;          // mm_interconnect_0:io_bridge_1_avalon_slave_0_write -> io_bridge_1:avs_write
	wire   [7:0] mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata;      // mm_interconnect_0:io_bridge_1_avalon_slave_0_writedata -> io_bridge_1:avs_writedata
	wire  [31:0] mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata;      // avalon2mem_0:avs_readdata -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest;   // avalon2mem_0:avs_waitrequest -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_waitrequest
	wire  [25:0] mm_interconnect_0_avalon2mem_0_avalon_slave_0_address;       // mm_interconnect_0:avalon2mem_0_avalon_slave_0_address -> avalon2mem_0:avs_address
	wire         mm_interconnect_0_avalon2mem_0_avalon_slave_0_read;          // mm_interconnect_0:avalon2mem_0_avalon_slave_0_read -> avalon2mem_0:avs_read
	wire   [3:0] mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable;    // mm_interconnect_0:avalon2mem_0_avalon_slave_0_byteenable -> avalon2mem_0:avs_byteenable
	wire         mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid; // avalon2mem_0:avs_readdatavalid -> mm_interconnect_0:avalon2mem_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_avalon2mem_0_avalon_slave_0_write;         // mm_interconnect_0:avalon2mem_0_avalon_slave_0_write -> avalon2mem_0:avs_write
	wire  [31:0] mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata;     // mm_interconnect_0:avalon2mem_0_avalon_slave_0_writedata -> avalon2mem_0:avs_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [8:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // io_bridge_0:avs_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // io_bridge_1:avs_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [avalon2mem_0:reset, io_bridge_0:reset, io_bridge_1:reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	avalon_to_mem32_bridge #(
		.g_tag (8'b01011011)
	) avalon2mem_0 (
		.reset               (rst_controller_reset_out_reset),                              //          reset.reset
		.avs_read            (mm_interconnect_0_avalon2mem_0_avalon_slave_0_read),          // avalon_slave_0.read
		.avs_write           (mm_interconnect_0_avalon2mem_0_avalon_slave_0_write),         //               .write
		.avs_address         (mm_interconnect_0_avalon2mem_0_avalon_slave_0_address),       //               .address
		.avs_writedata       (mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata),     //               .writedata
		.avs_byteenable      (mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable),    //               .byteenable
		.avs_waitrequest     (mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest),   //               .waitrequest
		.avs_readdata        (mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata),      //               .readdata
		.avs_readdatavalid   (mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid), //               .readdatavalid
		.clock               (clk_clk),                                                     //          clock.clk
		.mem_req_address     (mem_mem_req_address),                                         //            mem.mem_req_address
		.mem_req_byte_en     (mem_mem_req_byte_en),                                         //               .mem_req_byte_en
		.mem_req_read_writen (mem_mem_req_read_writen),                                     //               .mem_req_read_writen
		.mem_req_request     (mem_mem_req_request),                                         //               .mem_req_request
		.mem_req_tag         (mem_mem_req_tag),                                             //               .mem_req_tag
		.mem_req_wdata       (mem_mem_req_wdata),                                           //               .mem_req_wdata
		.mem_resp_dack_tag   (mem_mem_resp_dack_tag),                                       //               .mem_resp_dack_tag
		.mem_resp_data       (mem_mem_resp_data),                                           //               .mem_resp_data
		.mem_resp_rack_tag   (mem_mem_resp_rack_tag)                                        //               .mem_resp_rack_tag
	);

	avalon_to_io_bridge io_bridge_0 (
		.reset             (rst_controller_reset_out_reset),                             //          reset.reset
		.avs_read          (mm_interconnect_0_io_bridge_0_avalon_slave_0_read),          // avalon_slave_0.read
		.avs_write         (mm_interconnect_0_io_bridge_0_avalon_slave_0_write),         //               .write
		.avs_address       (mm_interconnect_0_io_bridge_0_avalon_slave_0_address),       //               .address
		.avs_writedata     (mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata),     //               .writedata
		.avs_ready         (mm_interconnect_0_io_bridge_0_avalon_slave_0_waitrequest),   //               .waitrequest_n
		.avs_readdata      (mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata),      //               .readdata
		.avs_readdatavalid (mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid), //               .readdatavalid
		.clock             (clk_clk),                                                    //          clock.clk
		.io_ack            (io_ack),                                                     //             io.ack
		.io_rdata          (io_rdata),                                                   //               .rdata
		.io_read           (io_read),                                                    //               .read
		.io_wdata          (io_wdata),                                                   //               .wdata
		.io_write          (io_write),                                                   //               .write
		.io_address        (io_address),                                                 //               .address
		.io_irq            (io_irq),                                                     //               .irq
		.avs_irq           (irq_mapper_receiver0_irq)                                    //            irq.irq
	);

	avalon_to_io_bridge io_bridge_1 (
		.reset             (rst_controller_reset_out_reset),                             //          reset.reset
		.avs_read          (mm_interconnect_0_io_bridge_1_avalon_slave_0_read),          // avalon_slave_0.read
		.avs_write         (mm_interconnect_0_io_bridge_1_avalon_slave_0_write),         //               .write
		.avs_address       (mm_interconnect_0_io_bridge_1_avalon_slave_0_address),       //               .address
		.avs_writedata     (mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata),     //               .writedata
		.avs_ready         (mm_interconnect_0_io_bridge_1_avalon_slave_0_waitrequest),   //               .waitrequest_n
		.avs_readdata      (mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata),      //               .readdata
		.avs_readdatavalid (mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid), //               .readdatavalid
		.clock             (clk_clk),                                                    //          clock.clk
		.io_ack            (io_u2p_ack),                                                 //             io.ack
		.io_rdata          (io_u2p_rdata),                                               //               .rdata
		.io_read           (io_u2p_read),                                                //               .read
		.io_wdata          (io_u2p_wdata),                                               //               .wdata
		.io_write          (io_u2p_write),                                               //               .write
		.io_address        (io_u2p_address),                                             //               .address
		.io_irq            (io_u2p_irq),                                                 //               .irq
		.avs_irq           (irq_mapper_receiver1_irq)                                    //            irq.irq
	);

	nios_solo_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_solo_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_solo_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.avalon2mem_0_avalon_slave_0_address            (mm_interconnect_0_avalon2mem_0_avalon_slave_0_address),       //              avalon2mem_0_avalon_slave_0.address
		.avalon2mem_0_avalon_slave_0_write              (mm_interconnect_0_avalon2mem_0_avalon_slave_0_write),         //                                         .write
		.avalon2mem_0_avalon_slave_0_read               (mm_interconnect_0_avalon2mem_0_avalon_slave_0_read),          //                                         .read
		.avalon2mem_0_avalon_slave_0_readdata           (mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdata),      //                                         .readdata
		.avalon2mem_0_avalon_slave_0_writedata          (mm_interconnect_0_avalon2mem_0_avalon_slave_0_writedata),     //                                         .writedata
		.avalon2mem_0_avalon_slave_0_byteenable         (mm_interconnect_0_avalon2mem_0_avalon_slave_0_byteenable),    //                                         .byteenable
		.avalon2mem_0_avalon_slave_0_readdatavalid      (mm_interconnect_0_avalon2mem_0_avalon_slave_0_readdatavalid), //                                         .readdatavalid
		.avalon2mem_0_avalon_slave_0_waitrequest        (mm_interconnect_0_avalon2mem_0_avalon_slave_0_waitrequest),   //                                         .waitrequest
		.io_bridge_0_avalon_slave_0_address             (mm_interconnect_0_io_bridge_0_avalon_slave_0_address),        //               io_bridge_0_avalon_slave_0.address
		.io_bridge_0_avalon_slave_0_write               (mm_interconnect_0_io_bridge_0_avalon_slave_0_write),          //                                         .write
		.io_bridge_0_avalon_slave_0_read                (mm_interconnect_0_io_bridge_0_avalon_slave_0_read),           //                                         .read
		.io_bridge_0_avalon_slave_0_readdata            (mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata),       //                                         .readdata
		.io_bridge_0_avalon_slave_0_writedata           (mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata),      //                                         .writedata
		.io_bridge_0_avalon_slave_0_readdatavalid       (mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid),  //                                         .readdatavalid
		.io_bridge_0_avalon_slave_0_waitrequest         (~mm_interconnect_0_io_bridge_0_avalon_slave_0_waitrequest),   //                                         .waitrequest
		.io_bridge_1_avalon_slave_0_address             (mm_interconnect_0_io_bridge_1_avalon_slave_0_address),        //               io_bridge_1_avalon_slave_0.address
		.io_bridge_1_avalon_slave_0_write               (mm_interconnect_0_io_bridge_1_avalon_slave_0_write),          //                                         .write
		.io_bridge_1_avalon_slave_0_read                (mm_interconnect_0_io_bridge_1_avalon_slave_0_read),           //                                         .read
		.io_bridge_1_avalon_slave_0_readdata            (mm_interconnect_0_io_bridge_1_avalon_slave_0_readdata),       //                                         .readdata
		.io_bridge_1_avalon_slave_0_writedata           (mm_interconnect_0_io_bridge_1_avalon_slave_0_writedata),      //                                         .writedata
		.io_bridge_1_avalon_slave_0_readdatavalid       (mm_interconnect_0_io_bridge_1_avalon_slave_0_readdatavalid),  //                                         .readdatavalid
		.io_bridge_1_avalon_slave_0_waitrequest         (~mm_interconnect_0_io_bridge_1_avalon_slave_0_waitrequest),   //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken)                  //                                         .clken
	);

	nios_solo_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
