library ieee;
use ieee.std_logic_1164.all;

package rocket_pkg is

    type t_byte_array is array (natural range <>) of std_logic_vector(7 downto 0);

    constant rocket_array : t_byte_array(0 to 7144) := (
        X"01", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"2D", X"31", X"7F", X"BF", X"7F", 
        X"BF", X"7F", X"EB", X"6A", X"EA", X"49", X"AC", X"B6", X"C9", X"6B", X"6B", X"A9", X"AA", X"B6", X"C9", X"AA", 
        X"EA", X"AB", X"2C", X"EA", X"C9", X"6D", X"6B", X"C9", X"AC", X"F6", X"C9", X"6B", X"6B", X"AA", X"EC", X"EA", 
        X"CF", X"26", X"9E", X"C9", X"2D", X"AB", X"A9", X"AC", X"B6", X"CB", X"6A", X"9A", X"49", X"AC", X"AA", X"A9", 
        X"2D", X"6B", X"69", X"ED", X"9A", X"6F", X"26", X"9E", X"C9", X"2D", X"9B", X"6B", X"6C", X"B5", X"AD", X"A7", 
        X"72", X"C9", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"64", X"92", X"49", X"64", X"92", X"4D", X"34", X"D6", X"49", X"B5", X"52", X"D9", X"37", X"95", X"AB", X"26", 
        X"93", X"4D", X"66", X"D3", X"5B", X"2C", X"9D", X"6D", X"B4", X"B2", X"AD", X"B5", X"B6", X"C9", X"67", X"53", 
        X"55", X"6D", X"9B", X"4A", X"D6", X"F3", X"69", X"A5", X"B2", X"C9", X"67", X"53", X"49", X"65", X"93", X"59", 
        X"35", X"52", X"B5", X"34", X"B3", X"AB", X"26", X"93", X"59", X"55", X"9D", X"55", X"2D", X"56", X"A9", X"A7", 
        X"73", X"6B", X"26", X"93", X"4D", X"65", X"75", X"A9", X"A4", X"B6", X"AD", X"34", X"D5", X"49", X"B5", X"52", 
        X"C9", X"27", X"9E", X"4F", X"37", X"B6", X"49", X"B5", X"B2", X"C9", X"27", X"96", X"4D", X"BC", X"96", X"4F", 
        X"57", X"76", X"6A", X"B6", X"B3", X"D5", X"54", X"D5", X"C9", X"24", X"F6", X"49", X"25", X"92", X"AD", X"35", 
        X"B6", X"57", X"27", X"95", X"69", X"64", X"D2", X"69", X"37", X"B2", X"5A", X"B6", X"93", X"A9", X"24", X"92", 
        X"A9", X"37", X"B2", X"5A", X"B6", X"D3", X"A9", X"64", X"D2", X"BB", X"2B", X"9A", X"55", X"ED", X"92", X"D7", 
        X"66", X"B5", X"59", X"5D", X"5B", X"4D", X"3C", X"9E", X"BB", X"6C", X"DD", X"4D", X"AB", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4A", X"AB", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"5F", X"EB", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", 
        X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"4B", X"46", X"E9", X"AA", X"FF", X"EB", 
        X"C9", X"2B", X"B6", X"4B", X"7F", X"EA", X"FF", X"EA", X"49", X"AC", X"B6", X"C9", X"7F", X"EB", X"7F", X"EB", 
        X"A9", X"AA", X"B6", X"C9", X"AA", X"FF", X"EA", X"AB", X"2C", X"FF", X"EA", X"C9", X"7F", X"ED", X"7F", X"EB", 
        X"C9", X"AC", X"F6", X"C9", X"7F", X"EB", X"7F", X"EB", X"AA", X"FF", X"EC", X"FF", X"EA", X"CF", X"26", X"9E", 
        X"C9", X"2D", X"AB", X"A9", X"AC", X"B6", X"CB", X"7F", X"EA", X"9A", X"49", X"AC", X"AA", X"A9", X"2D", X"7F", 
        X"EB", X"7F", X"E9", X"FF", X"ED", X"9A", X"7F", X"EF", X"26", X"9E", X"C9", X"2D", X"9B", X"7F", X"EB", X"7F", 
        X"EC", X"B5", X"AD", X"A7", X"72", X"C9", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"7F", X"E4", X"92", X"49", X"7F", X"E4", X"92", X"4D", X"34", X"D6", X"49", X"B5", 
        X"52", X"D9", X"37", X"95", X"AB", X"26", X"93", X"4D", X"7F", X"E6", X"D3", X"5B", X"2C", X"9D", X"7F", X"ED", 
        X"B4", X"B2", X"AD", X"B5", X"B6", X"C9", X"7F", X"E7", X"53", X"55", X"7F", X"ED", X"9B", X"4A", X"D6", X"F3", 
        X"7F", X"E9", X"A5", X"B2", X"C9", X"7F", X"E7", X"53", X"49", X"7F", X"E5", X"93", X"59", X"35", X"52", X"B5", 
        X"34", X"B3", X"AB", X"26", X"93", X"59", X"55", X"9D", X"55", X"2D", X"56", X"A9", X"A7", X"73", X"7F", X"EB", 
        X"26", X"93", X"4D", X"7F", X"E5", X"75", X"A9", X"A4", X"B6", X"AD", X"34", X"D5", X"49", X"B5", X"52", X"C9", 
        X"27", X"9E", X"4F", X"37", X"B6", X"49", X"B5", X"B2", X"C9", X"27", X"96", X"4D", X"BC", X"96", X"4F", X"57", 
        X"76", X"7F", X"EA", X"B6", X"B3", X"D5", X"54", X"D5", X"C9", X"24", X"F6", X"49", X"25", X"92", X"AD", X"35", 
        X"B6", X"57", X"27", X"95", X"7F", X"E9", X"7F", X"E4", X"D2", X"7F", X"E9", X"37", X"B2", X"5A", X"B6", X"93", 
        X"A9", X"24", X"92", X"A9", X"37", X"B2", X"5A", X"B6", X"D3", X"A9", X"7F", X"E4", X"D2", X"BB", X"2B", X"9A", 
        X"55", X"FF", X"ED", X"92", X"D7", X"7F", X"E6", X"B5", X"59", X"5D", X"5B", X"4D", X"3C", X"9E", X"BB", X"7F", 
        X"EC", X"DD", X"4D", X"A5", X"96", X"CB", X"25", X"96", X"55", X"2B", X"72", X"49", X"24", X"9B", X"D9", X"5D", 
        X"AD", X"7F", X"ED", X"24", X"9D", X"4B", X"7F", X"EA", X"FF", X"EA", X"C9", X"FF", X"EC", X"FF", X"EB", X"4E", 
        X"A6", X"FF", X"EE", X"4F", X"26", X"9D", X"7F", X"EA", X"AB", X"7F", X"EA", X"7F", X"ED", X"7F", X"E4", X"DE", 
        X"AA", X"AB", X"7F", X"EA", X"4D", X"7F", X"E4", X"DE", X"4A", X"AA", X"AA", X"49", X"AA", X"9A", X"7F", X"E9", 
        X"2A", X"D6", X"49", X"AA", X"9B", X"C9", X"7F", X"ED", X"7F", X"EB", X"CA", X"FF", X"EA", X"AA", X"AF", X"26", 
        X"9E", X"C9", X"AD", X"76", X"C9", X"FF", X"EC", X"DB", X"7F", X"ED", X"24", X"9D", X"AB", X"2B", X"AA", X"C9", 
        X"2C", X"FF", X"EB", X"4D", X"A7", X"72", X"C9", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"4D", X"59", X"29", X"24", X"92", X"49", X"24", X"96", X"49", X"BA", 
        X"F2", X"57", X"7F", X"E7", X"76", X"49", X"D4", X"F2", X"4D", X"35", X"B6", X"49", X"B5", X"B2", X"D9", X"37", 
        X"95", X"79", X"34", X"B2", X"B9", X"B5", X"95", X"A9", X"24", X"FF", X"EB", X"4F", X"57", X"73", X"49", X"2D", 
        X"9B", X"C9", X"25", X"92", X"AD", X"7F", X"E4", X"DE", X"7F", X"EA", X"AB", X"7F", X"EA", X"CB", X"7F", X"ED", 
        X"7F", X"EA", X"49", X"7F", X"ED", X"7F", X"EA", X"AB", X"2B", X"9A", X"CF", X"26", X"92", X"7F", X"EF", X"25", 
        X"B3", X"4D", X"A6", X"F2", X"C9", X"2D", X"9A", X"7F", X"E9", X"2A", X"DA", X"7F", X"E9", X"AD", X"9A", X"4F", 
        X"7F", X"E6", X"DE", X"7F", X"E9", X"AC", X"AA", X"7F", X"E9", X"AD", X"9A", X"7F", X"E9", X"2B", X"B6", X"4D", 
        X"24", X"9E", X"7F", X"E9", X"AD", X"9B", X"4F", X"7F", X"E6", X"DE", X"49", X"7F", X"ED", X"7F", X"EA", X"AB", 
        X"2B", X"9A", X"C9", X"2A", X"F6", X"49", X"2A", X"DA", X"A9", X"2A", X"FF", X"EA", X"AB", X"7F", X"EC", X"9A", 
        X"C9", X"AC", X"AA", X"4D", X"A5", X"52", X"CD", X"24", X"96", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", 
        X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"55", X"95", 
        X"2F", X"26", X"9A", X"D9", X"34", X"B6", X"59", X"34", X"93", X"5B", X"2C", X"9D", X"AD", X"7F", X"E4", X"DE", 
        X"D9", X"34", X"B2", X"A9", X"25", X"95", X"75", X"B7", X"76", X"7B", X"35", X"9E", X"55", X"BD", X"AD", X"B7", 
        X"37", X"B2", X"4D", X"A4", X"92", X"C9", X"AC", X"D2", X"A9", X"B4", X"B3", X"AF", X"7F", X"E7", X"73", X"AA", 
        X"B6", X"B3", X"AD", X"A4", X"95", X"C9", X"2A", X"92", X"AD", X"7F", X"E4", X"DE", X"D9", X"34", X"B2", X"B9", 
        X"BC", X"95", X"B9", X"34", X"D3", X"AB", X"26", X"93", X"57", X"56", X"DE", X"A9", X"A4", X"96", X"4B", X"27", 
        X"B2", X"49", X"24", X"FF", X"EB", X"C9", X"A7", X"92", X"75", X"54", X"DB", X"59", X"34", X"F5", X"AB", X"26", 
        X"93", X"D7", X"57", X"7F", X"EA", X"C9", X"B5", X"B2", X"D9", X"B7", X"96", X"D9", X"34", X"93", X"CB", X"26", 
        X"93", X"4D", X"B5", X"B6", X"CB", X"25", X"96", X"57", X"34", X"9E", X"4D", X"BA", X"92", X"C9", X"25", X"92", 
        X"AF", X"37", X"B6", X"C9", X"D4", X"FF", X"EA", X"4D", X"35", X"B6", X"7F", X"ED", X"A5", X"96", X"DB", X"35", 
        X"9A", X"4F", X"36", X"F2", X"59", X"D7", X"9B", X"DB", X"7F", X"EC", X"DE", X"DB", X"27", X"9A", X"55", X"7F", 
        X"EA", X"AE", X"DA", X"BA", X"DA", X"D5", X"AD", X"7F", X"EE", X"57", X"36", X"9A", X"55", X"2D", X"B6", X"D5", 
        X"34", X"93", X"79", X"36", X"D2", X"A9", X"27", X"96", X"49", X"D5", X"92", X"AD", X"55", X"7F", X"EE", X"49", 
        X"B5", X"B2", X"DA", X"B5", X"9A", X"C9", X"3B", X"AB", X"CD", X"2B", X"56", X"7F", X"ED", X"35", X"92", X"CB", 
        X"27", X"92", X"49", X"A4", X"D6", X"CD", X"36", X"96", X"A9", X"AD", X"92", X"C9", X"A4", X"FF", X"EB", X"4D", 
        X"2B", X"56", X"7F", X"EE", X"B6", X"B5", X"CD", X"34", X"D6", X"7F", X"E9", X"DC", X"F6", X"CF", X"3C", X"93", 
        X"4D", X"DC", X"F2", X"C9", X"26", X"92", X"DB", X"5B", X"7F", X"ED", X"B7", X"7F", X"E6", X"9B", X"B9", X"35", 
        X"55", X"55", X"25", X"B2", X"49", X"D4", X"FF", X"EA", X"4B", X"37", X"53", X"4D", X"AD", X"B6", X"C9", X"A7", 
        X"95", X"B9", X"34", X"F2", X"B5", X"34", X"B3", X"AB", X"26", X"93", X"D7", X"37", X"AB", X"C9", X"A4", X"B6", 
        X"A9", X"B5", X"B2", X"D9", X"B7", X"96", X"79", X"BC", X"D3", X"CF", X"5C", X"D6", X"49", X"B5", X"B2", X"79", 
        X"37", X"95", X"AA", X"A6", X"B3", X"D7", X"54", X"DB", X"7F", X"ED", X"D4", X"FF", X"EE", X"49", X"DC", X"F2", 
        X"57", X"7F", X"EC", X"DD", X"49", X"DC", X"9A", X"5B", X"7F", X"EC", X"DA", X"CE", X"B6", X"B5", X"C9", X"D4", 
        X"F6", X"CD", X"34", X"D6", X"7F", X"EB", X"5B", X"72", X"4D", X"36", X"96", X"7B", X"2B", X"55", X"AD", X"56", 
        X"D6", X"C9", X"D4", X"FF", X"EA", X"AD", X"B5", X"B6", X"C9", X"A7", X"95", X"AA", X"B5", X"53", X"7F", X"ED", 
        X"54", X"D6", X"C9", X"B5", X"B2", X"C9", X"A7", X"9E", X"CD", X"B5", X"B6", X"DA", X"B6", X"DA", X"C9", X"24", 
        X"F6", X"49", X"3D", X"72", X"B5", X"54", X"D5", X"D9", X"34", X"F5", X"79", X"35", X"92", X"AD", X"2D", X"52", 
        X"49", X"2A", X"92", X"CD", X"A4", X"95", X"C9", X"7F", X"E6", X"D2", X"54", X"BC", X"B6", X"A6", X"AA", X"7F", 
        X"E9", X"3D", X"B2", X"4D", X"3A", X"96", X"A9", X"DC", X"9D", X"D9", X"7F", X"EA", X"DD", X"AD", X"2C", X"92", 
        X"4D", X"AA", X"96", X"AD", X"35", X"B6", X"75", X"25", X"53", X"4D", X"A5", X"96", X"CB", X"25", X"96", X"5B", 
        X"37", X"7F", X"EA", X"59", X"B5", X"9B", X"DB", X"7F", X"EC", X"DE", X"D7", X"2B", X"9E", X"55", X"2A", X"F5", 
        X"CB", X"26", X"93", X"4A", X"FF", X"EB", X"5D", X"C9", X"24", X"B6", X"CB", X"27", X"9E", X"49", X"A4", X"F6", 
        X"C9", X"7F", X"E4", X"D2", X"55", X"7F", X"EA", X"DE", X"B9", X"7F", X"EA", X"DA", X"57", X"36", X"9B", X"B9", 
        X"D4", X"9A", X"5A", X"BA", X"9E", X"D5", X"26", X"D2", X"AB", X"25", X"B3", X"4D", X"2D", X"B6", X"C9", X"DC", 
        X"FF", X"EA", X"A9", X"56", X"D2", X"4D", X"DC", X"FF", X"EE", X"AA", X"B6", X"B3", X"B9", X"7F", X"EA", X"D5", 
        X"AE", X"BA", X"D5", X"CE", X"B6", X"D5", X"CD", X"3C", X"93", X"79", X"26", X"96", X"D7", X"24", X"95", X"75", 
        X"7F", X"E5", X"7F", X"EB", X"C9", X"B5", X"B3", X"59", X"B7", X"95", X"AA", X"AB", X"5A", X"D6", X"AD", X"53", 
        X"C9", X"AD", X"B2", X"BA", X"B5", X"9A", X"CE", X"BC", X"DE", X"D6", X"AD", X"53", X"CD", X"B5", X"B6", X"AA", 
        X"A5", X"96", X"CB", X"27", X"9A", X"56", X"AD", X"53", X"CD", X"B5", X"B6", X"AA", X"A5", X"92", X"CA", X"A7", 
        X"9A", X"D6", X"AD", X"53", X"C9", X"AD", X"B2", X"B9", X"B7", X"9A", X"7B", X"35", X"AA", X"5A", X"AD", X"9E", 
        X"D5", X"AD", X"9D", X"B6", X"BA", X"9E", X"D9", X"AA", X"D6", X"D9", X"34", X"92", X"CF", X"25", X"5E", X"56", 
        X"AD", X"53", X"CD", X"B5", X"56", X"BA", X"B5", X"95", X"CB", X"24", X"95", X"AD", X"B7", X"B6", X"CA", X"A6", 
        X"DA", X"CD", X"DB", X"95", X"D9", X"35", X"52", X"B9", X"DA", X"F5", X"4B", X"26", X"B3", X"C9", X"AB", X"B2", 
        X"DA", X"B6", X"D3", X"A9", X"7F", X"E4", X"D2", X"4A", X"FF", X"EA", X"F5", X"CA", X"D6", X"F5", X"CE", X"B6", 
        X"AE", X"7F", X"E9", X"7F", X"E5", X"93", X"4A", X"B6", X"AA", X"7F", X"ED", X"B5", X"56", X"AA", X"A5", X"9B", 
        X"7F", X"E9", X"7F", X"E4", X"D2", X"CB", X"35", X"AA", X"49", X"24", X"DA", X"B5", X"37", X"56", X"B5", X"37", 
        X"52", X"A9", X"FF", X"EA", X"F3", X"D9", X"55", X"95", X"CB", X"26", X"B3", X"C9", X"AB", X"B2", X"DA", X"B6", 
        X"D3", X"AD", X"54", X"D6", X"4A", X"FF", X"EA", X"F5", X"CA", X"D6", X"F5", X"DB", X"2B", X"9A", X"55", X"A7", 
        X"B3", X"B5", X"AD", X"95", X"7F", X"EA", X"A7", X"93", X"7F", X"EE", X"D6", X"F3", X"CB", X"3A", X"9A", X"4D", 
        X"5A", X"D6", X"57", X"7F", X"E7", X"7F", X"EB", X"B5", X"3C", X"92", X"5B", X"36", X"93", X"49", X"7F", X"ED", 
        X"9B", X"49", X"7F", X"ED", X"9B", X"49", X"37", X"B2", X"59", X"B4", X"F3", X"DB", X"2C", X"9E", X"AD", X"35", 
        X"B6", X"C9", X"A5", X"B2", X"D9", X"B7", X"9B", X"7F", X"EB", X"26", X"93", X"C9", X"25", X"93", X"79", X"35", 
        X"93", X"AB", X"26", X"93", X"D7", X"37", X"9A", X"59", X"B5", X"55", X"B5", X"7F", X"E4", X"D3", X"49", X"B5", 
        X"B2", X"7F", X"E9", X"27", X"95", X"CA", X"A6", X"B3", X"D7", X"54", X"DB", X"74", X"B5", X"AB", X"3B", X"56", 
        X"55", X"AA", X"B3", X"B5", X"34", X"96", X"AD", X"24", X"9A", X"4D", X"35", X"B6", X"57", X"27", X"95", X"7F", 
        X"E9", X"7F", X"E4", X"D2", X"5B", X"2B", X"9A", X"55", X"2B", X"53", X"79", X"25", X"93", X"AD", X"55", X"76", 
        X"57", X"27", X"B5", X"B9", X"FF", X"E5", X"75", X"C9", X"24", X"DE", X"4D", X"24", X"95", X"49", X"A4", X"B6", 
        X"C9", X"D5", X"92", X"AE", X"B6", X"B5", X"C9", X"D4", X"F3", X"4E", X"B6", X"B5", X"A9", X"D4", X"F3", X"7F", 
        X"ED", X"A4", X"95", X"AF", X"7F", X"EC", X"D3", X"AD", X"A4", X"95", X"CD", X"2A", X"93", X"55", X"54", X"D2", 
        X"C9", X"A4", X"B6", X"CD", X"37", X"56", X"AD", X"24", X"95", X"49", X"A4", X"B6", X"CD", X"B4", X"D6", X"7F", 
        X"ED", X"55", X"76", X"49", X"B5", X"B2", X"D9", X"37", X"95", X"7F", X"E9", X"36", X"96", X"49", X"36", X"92", 
        X"A9", X"56", X"D3", X"55", X"54", X"D5", X"59", X"B4", X"B5", X"A9", X"36", X"96", X"49", X"36", X"92", X"AD", 
        X"56", X"D6", X"7F", X"EF", X"26", X"9A", X"C9", X"24", X"AB", X"CD", X"7F", X"E7", X"B6", X"77", X"27", X"B2", 
        X"57", X"36", X"96", X"5A", X"B6", X"B2", X"CD", X"3A", X"F2", X"49", X"35", X"52", X"B7", X"27", X"B2", X"57", 
        X"36", X"96", X"5A", X"B6", X"B2", X"D7", X"2B", X"B2", X"55", X"2D", X"53", X"7F", X"E9", X"34", X"96", X"49", 
        X"36", X"92", X"A9", X"56", X"D3", X"CD", X"5C", X"D5", X"77", X"7F", X"EC", X"DD", X"B5", X"54", X"D5", X"59", 
        X"B4", X"B5", X"A9", X"34", X"96", X"49", X"36", X"92", X"B7", X"24", X"9E", X"AF", X"26", X"9A", X"C9", X"24", 
        X"B6", X"4D", X"37", X"56", X"B9", X"2A", X"9B", X"AD", X"34", X"96", X"75", X"25", X"AE", X"49", X"5A", X"D2", 
        X"4D", X"34", X"96", X"B9", X"3B", X"92", X"B9", X"D4", X"D6", X"4A", X"A6", X"96", X"D5", X"AB", X"9A", X"CB", 
        X"26", X"B3", X"4D", X"3A", X"96", X"DB", X"27", X"9A", X"4F", X"3C", X"B3", X"55", X"3B", X"92", X"49", X"24", 
        X"9E", X"4F", X"26", X"9A", X"D9", X"34", X"B5", X"7F", X"E9", X"24", X"B5", X"CB", X"26", X"93", X"57", X"7F", 
        X"EC", X"DB", X"7F", X"ED", X"7F", X"E4", X"DE", X"DB", X"36", X"B3", X"7F", X"E9", X"7F", X"E4", X"D2", X"BB", 
        X"2B", X"9A", X"4D", X"BA", X"FF", X"EA", X"D7", X"56", X"D3", X"A9", X"A4", X"D6", X"C9", X"BA", X"F2", X"4D", 
        X"B5", X"B6", X"DA", X"B6", X"DE", X"C9", X"24", X"F6", X"49", X"3D", X"72", X"B9", X"BD", X"9D", X"59", X"B4", 
        X"B5", X"7F", X"ED", X"BB", X"56", X"7F", X"EB", X"7F", X"EB", X"73", X"BA", X"FF", X"E7", X"7F", X"ED", X"59", 
        X"B4", X"B5", X"7F", X"E9", X"7F", X"E4", X"D2", X"C9", X"7F", X"ED", X"73", X"A9", X"B5", X"B2", X"D9", X"B4", 
        X"D5", X"7F", X"ED", X"FF", X"E5", X"96", X"49", X"2D", X"B3", X"C9", X"D5", X"75", X"59", X"B4", X"D5", X"7F", 
        X"E9", X"7F", X"ED", X"72", X"C9", X"7F", X"ED", X"73", X"A9", X"B5", X"AB", X"A9", X"A4", X"DE", X"CD", X"55", 
        X"76", X"49", X"B5", X"B2", X"D9", X"37", X"95", X"7F", X"E9", X"A4", X"95", X"4B", X"26", X"93", X"57", X"7F", 
        X"EC", X"DB", X"7F", X"ED", X"A5", X"96", X"DB", X"35", X"9A", X"55", X"2B", X"72", X"5B", X"5B", X"95", X"D6", 
        X"93", X"29", X"FF", X"E5", X"B2", X"CD", X"B7", X"B6", X"C9", X"A4", X"FF", X"EB", X"C9", X"35", X"55", X"79", 
        X"D5", X"B6", X"D9", X"54", X"D3", X"CB", X"26", X"93", X"4D", X"B5", X"56", X"DB", X"35", X"9E", X"55", X"7F", 
        X"EB", X"B3", X"CB", X"26", X"93", X"49", X"3A", X"92", X"49", X"3A", X"92", X"49", X"B5", X"B2", X"C9", X"7F", 
        X"E7", X"53", X"4D", X"7F", X"E5", X"75", X"49", X"B5", X"B2", X"C9", X"27", X"9D", X"49", X"B5", X"B2", X"C9", 
        X"7F", X"E7", X"53", X"4D", X"7F", X"E5", X"75", X"49", X"B5", X"B2", X"DB", X"35", X"95", X"7F", X"E9", X"7F", 
        X"EB", X"92", X"4D", X"35", X"53", X"79", X"B5", X"73", X"7F", X"EB", X"26", X"93", X"49", X"25", X"55", X"79", 
        X"35", X"53", X"AB", X"26", X"93", X"4D", X"B7", X"B6", X"D9", X"B4", X"F3", X"7F", X"EB", X"26", X"93", X"49", 
        X"25", X"55", X"79", X"35", X"53", X"AB", X"26", X"93", X"55", X"27", X"B2", X"B9", X"54", X"95", X"4D", X"7F", 
        X"E5", X"75", X"A9", X"B5", X"B2", X"C9", X"7F", X"E7", X"53", X"4D", X"7F", X"E5", X"75", X"49", X"B5", X"B2", 
        X"DB", X"35", X"95", X"A9", X"7F", X"E4", X"D2", X"A9", X"B5", X"B2", X"C9", X"7F", X"E7", X"53", X"4D", X"7F", 
        X"E5", X"75", X"49", X"B5", X"B2", X"D9", X"37", X"93", X"5B", X"34", X"93", X"7F", X"ED", X"55", X"76", X"49", 
        X"B5", X"B2", X"C9", X"27", X"9E", X"55", X"7F", X"E7", X"AE", X"55", X"7F", X"E6", X"FF", X"EE", X"56", X"FF", 
        X"E4", X"B3", X"7F", X"EF", X"7F", X"EC", X"9A", X"7F", X"EE", X"AC", X"9A", X"7F", X"EE", X"FF", X"EC", X"9A", 
        X"7F", X"EF", X"2D", X"9B", X"7F", X"EF", X"7F", X"ED", X"9B", X"7F", X"EE", X"AD", X"9B", X"7F", X"EE", X"FF", 
        X"ED", X"9B", X"79", X"24", X"92", X"79", X"7F", X"E4", X"92", X"79", X"A4", X"92", X"79", X"FF", X"E4", X"92", 
        X"79", X"25", X"93", X"79", X"7F", X"E5", X"93", X"79", X"A5", X"93", X"79", X"FF", X"E5", X"93", X"7B", X"24", 
        X"92", X"7F", X"EF", X"7F", X"E5", X"B3", X"4F", X"25", X"B3", X"4E", X"A5", X"92", X"7F", X"EE", X"A4", X"F3", 
        X"AF", X"25", X"92", X"CF", X"7F", X"E5", X"52", X"7F", X"EF", X"24", X"D2", X"7F", X"ED", X"2D", X"9D", X"49", 
        X"24", X"95", X"CE", X"FF", X"E5", X"93", X"7F", X"EE", X"A5", X"B2", X"CB", X"7F", X"E6", X"D6", X"AD", X"FF", 
        X"E6", X"93", X"7F", X"ED", X"A5", X"53", X"4D", X"FF", X"E5", X"73", X"AA", X"FF", X"E4", X"F2", X"AD", X"24", 
        X"D6", X"4D", X"FF", X"E4", X"F3", X"CD", X"25", X"93", X"7F", X"E9", X"24", X"96", X"CD", X"FF", X"E4", X"B2", 
        X"4D", X"7F", X"E4", X"F2", X"77", X"36", X"93", X"7F", X"E9", X"7F", X"E4", X"D2", X"A9", X"37", X"B2", X"59", 
        X"34", X"D3", X"5B", X"7F", X"EC", X"DE", X"AF", X"7F", X"EA", X"D5", X"AA", X"A5", X"53", X"7F", X"EB", X"25", 
        X"73", X"CB", X"25", X"53", X"7F", X"EA", X"FF", X"E4", X"B3", X"4A", X"FF", X"E7", X"72", X"4A", X"FF", X"E5", 
        X"92", X"AB", X"7F", X"E5", X"B2", X"AB", X"26", X"92", X"CB", X"26", X"92", X"AB", X"7F", X"E4", X"92", X"7F", 
        X"EB", X"24", X"B3", X"49", X"FF", X"E5", X"B3", X"49", X"25", X"52", X"4A", X"A7", X"72", X"C9", X"A5", X"53", 
        X"7F", X"E9", X"25", X"53", X"C9", X"7F", X"E5", X"93", X"7F", X"E9", X"25", X"93", X"7F", X"E9", X"FF", X"E4", 
        X"B2", X"49", X"FF", X"E4", X"D2", X"49", X"A4", X"B2", X"49", X"7F", X"E4", X"92", X"7F", X"E9", X"24", X"B2", 
        X"4D", X"A5", X"93", X"49", X"AD", X"93", X"C9", X"A4", X"AB", X"4D", X"BD", X"96", X"7F", X"EE", X"99", X"2D", 
        X"34", X"96", X"4A", X"B6", X"96", X"CD", X"35", X"AA", X"5A", X"FF", X"E7", X"7F", X"ED", X"7F", X"E9", X"A4", 
        X"F6", X"CD", X"DB", X"B6", X"77", X"25", X"53", X"A9", X"24", X"92", X"7F", X"EA", X"B6", X"B6", X"AF", X"34", 
        X"B2", X"49", X"37", X"B2", X"59", X"B4", X"FF", X"EB", X"DB", X"2C", X"9D", X"4A", X"AB", X"93", X"7F", X"EA", 
        X"A6", X"FF", X"ED", X"CD", X"DC", X"92", X"CD", X"DC", X"92", X"D5", X"7F", X"E5", X"7F", X"EB", X"C9", X"B5", 
        X"B3", X"59", X"D7", X"56", X"D9", X"B4", X"B5", X"B9", X"AC", X"D3", X"7F", X"EB", X"26", X"93", X"D5", X"25", 
        X"B2", X"49", X"B5", X"B2", X"7F", X"E9", X"27", X"95", X"CA", X"A6", X"B3", X"D7", X"54", X"DB", X"75", X"37", 
        X"93", X"AB", X"26", X"93", X"CD", X"25", X"53", X"7F", X"E9", X"24", X"FF", X"EB", X"AB", X"26", X"93", X"DB", 
        X"2B", X"5A", X"55", X"AC", X"D2", X"D9", X"34", X"92", X"D5", X"B7", X"53", X"B9", X"34", X"B2", X"B5", X"36", 
        X"B3", X"79", X"34", X"F2", X"BB", X"36", X"95", X"5B", X"5C", X"DD", X"CD", X"B5", X"B6", X"B9", X"B7", X"9B", 
        X"BB", X"3D", X"5E", X"59", X"55", X"9B", X"5B", X"7F", X"EC", X"DE", X"7F", X"E9", X"BC", X"D2", X"D9", X"7F", 
        X"EA", X"DD", X"B9", X"BD", X"9B", X"B9", X"B4", X"F6", X"DB", X"36", X"D5", X"5B", X"5C", X"DD", X"CD", X"B5", 
        X"B6", X"B9", X"B7", X"9B", X"BB", X"3D", X"5E", X"56", X"AC", X"DD", X"AD", X"DC", X"96", X"7B", X"7F", X"EC", 
        X"DB", X"7F", X"EB", X"37", X"92", X"56", X"AB", X"53", X"CD", X"34", X"96", X"4A", X"D6", X"D5", X"DB", X"5C", 
        X"DD", X"D5", X"27", X"93", X"AB", X"26", X"B3", X"D7", X"57", X"72", X"C9", X"B4", X"B6", X"BB", X"5C", X"DD", 
        X"D5", X"27", X"93", X"AB", X"26", X"B3", X"D7", X"57", X"7F", X"ED", X"7F", X"E9", X"AC", X"B6", X"AB", X"34", 
        X"B6", X"4A", X"FF", X"EA", X"F5", X"CA", X"D6", X"F5", X"CB", X"3B", X"9A", X"56", X"AD", X"53", X"CD", X"B5", 
        X"B6", X"A9", X"A7", X"95", X"AD", X"AD", X"AE", X"77", X"36", X"B6", X"7F", X"ED", X"26", X"9E", X"B5", X"37", 
        X"56", X"B5", X"37", X"5D", X"5B", X"2C", X"9A", X"4D", X"54", X"96", X"5B", X"5C", X"DD", X"C9", X"AD", X"B2", 
        X"BA", X"B5", X"95", X"DB", X"2B", X"5A", X"55", X"AA", X"F3", X"CD", X"5A", X"D5", X"AD", X"35", X"B2", X"49", 
        X"B4", X"B6", X"D5", X"25", X"AB", X"C9", X"B5", X"B3", X"59", X"B7", X"B5", X"B5", X"3B", X"55", X"AB", X"26", 
        X"D3", X"55", X"3C", X"93", X"7F", X"E9", X"2D", X"9B", X"AB", X"26", X"93", X"C9", X"B5", X"B2", X"D9", X"B7", 
        X"95", X"B5", X"24", X"95", X"AA", X"A6", X"B3", X"CD", X"A5", X"96", X"7F", X"EB", X"25", X"96", X"55", X"2B", 
        X"73", X"AB", X"26", X"93", X"C9", X"2D", X"AB", X"49", X"B5", X"B2", X"C9", X"A7", X"9B", X"49", X"7F", X"ED", 
        X"72", X"B6", X"D4", X"AB", X"7F", X"E9", X"AA", X"B2", X"C9", X"24", X"92", X"49", X"24", X"92", X"49", X"24", 
        X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", 
        X"49", X"24", X"92", X"49", X"24", X"92", X"49", X"24", X"92", X"4D", X"29", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", X"69", 
        X"68", X"D6", X"96", X"96", X"96", X"96", X"96", X"96", X"96" );

end;
