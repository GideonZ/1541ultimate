
library ieee;
use ieee.std_logic_1164.all;

package bootrom_pkg is
    type t_boot_data    is array(natural range <>) of std_logic_vector(31 downto 0);

    constant c_bootrom : t_boot_data(0 to 2047) := (
        X"30047073", X"00002117", X"ff810113", X"00002197", X"3f418193", X"00000517", X"0cc50513", X"30551073",
        X"34151073", X"30001073", X"30401073", X"34401073", X"32001073", X"30601073", X"b0001073", X"b8001073",
        X"b0201073", X"b8201073", X"00000093", X"00000213", X"00000293", X"00000313", X"00000393", X"00001597",
        X"c7c58593", X"00002617", X"b9c60613", X"00002697", X"b9468693", X"00d65c63", X"0005a703", X"00e62023",
        X"00458593", X"00460613", X"fedff06f", X"00002717", X"b7470713", X"80818793", X"00f75863", X"00072023",
        X"00470713", X"ff5ff06f", X"00000513", X"00000593", X"088000ef", X"34051073", X"10500073", X"0000006f",
        X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013",
        X"ff810113", X"00812023", X"00912223", X"34202473", X"02044663", X"34102473", X"00041483", X"0034f493",
        X"00240413", X"34141073", X"00300413", X"00941863", X"34102473", X"00240413", X"34141073", X"10000437",
        X"04900493", X"00940fa3", X"00012403", X"00412483", X"00810113", X"30200073", X"fe010113", X"80001537",
        X"00812c23", X"01412423", X"10060437", X"00300a13", X"c0850513", X"00112e23", X"00912a23", X"01212823",
        X"01312623", X"01512223", X"fff00993", X"195000ef", X"21440423", X"21340023", X"00100a93", X"21540423",
        X"21340023", X"21440423", X"1d1000ef", X"00050493", X"10100937", X"3f8000ef", X"00c94503", X"0ff57513",
        X"17c000ef", X"0404d863", X"1c0000ef", X"1571c4b7", X"00010437", X"abe48493", X"800019b7", X"80001a37",
        X"ffc42783", X"14979663", X"c7498513", X"40c000ef", X"fe042e23", X"ff842903", X"00090513", X"3b0000ef",
        X"c48a0513", X"3f4000ef", X"00090513", X"12c000ef", X"fd1ff06f", X"70090423", X"478000ef", X"00010937",
        X"168000ef", X"ffc92703", X"1571c7b7", X"abe78793", X"02f71663", X"80001537", X"c2050513", X"3bc000ef",
        X"fe092e23", X"ff892503", X"0f0000ef", X"80001537", X"c4c50513", X"3a4000ef", X"f75ff06f", X"40000537",
        X"00a4f4b3", X"fe0494e3", X"21540423", X"21440023", X"02200793", X"20f40023", X"20040023", X"20040023",
        X"20042903", X"20042483", X"20042403", X"00090513", X"31c000ef", X"00048513", X"314000ef", X"00040513",
        X"30c000ef", X"80001537", X"c2850513", X"34c000ef", X"f9348ee3", X"001807b7", X"00090513", X"fff48493",
        X"ffe78793", X"10060737", X"0497f263", X"100607b7", X"80001537", X"20078423", X"c3850513", X"31c000ef",
        X"100007b7", X"00a7c783", X"0e07f793", X"01879793", X"4187d793", X"0207c663", X"00040513", X"03c000ef",
        X"00000013", X"00000013", X"ff9ff06f", X"20072683", X"ffc48493", X"00450513", X"fed52e23", X"fadff06f",
        X"80001537", X"c4450513", X"2d0000ef", X"fd5ff06f", X"00000013", X"eadff06f", X"00050067", X"ff010113",
        X"00812423", X"80001437", X"c7c40413", X"00455793", X"00f407b3", X"00912223", X"00050493", X"0007c503",
        X"00f4f493", X"00112623", X"00940433", X"075000ef", X"00044503", X"00812403", X"00c12083", X"00412483",
        X"01010113", X"05d0006f", X"050507b7", X"fe010113", X"05778793", X"00f12023", X"4a5357b7", X"4cf78793",
        X"00f12223", X"010107b7", X"05778793", X"00f12423", X"adcaa7b7", X"20f78793", X"00f12623", X"00112e23",
        X"00812c23", X"00912a23", X"10100437", X"70744503", X"0ff57513", X"f69ff0ef", X"00a00513", X"005000ef",
        X"00c44783", X"10100637", X"0ff7f793", X"0037d793", X"feb78793", X"00f03733", X"70e40323", X"fc800713",
        X"70e40023", X"70164703", X"01871713", X"41875713", X"14074663", X"01400713", X"70e60023", X"10100637",
        X"70164703", X"01871713", X"41875713", X"12074c63", X"00800713", X"70e60023", X"101006b7", X"7016c703",
        X"01871713", X"41875713", X"12074263", X"00000713", X"101005b7", X"00800513", X"00e106b3", X"0006c683",
        X"70d58023", X"7015c683", X"01869693", X"4186d693", X"1006c263", X"00170713", X"fea710e3", X"00100713",
        X"70e581a3", X"10100637", X"70164683", X"01869693", X"4186d693", X"0e06c463", X"0017b793", X"70f60323",
        X"fc800793", X"70f60023", X"101006b7", X"7016c783", X"01879793", X"4187d793", X"0c07c663", X"01400793",
        X"70f68023", X"101006b7", X"7016c783", X"01879793", X"4187d793", X"0a07cc63", X"00800793", X"70f68023",
        X"10100737", X"70174783", X"01879793", X"4187d793", X"0a07c263", X"00000793", X"10100637", X"00800593",
        X"00810713", X"00f70733", X"00074703", X"70e60023", X"70164703", X"01871713", X"41875713", X"08074063",
        X"00178793", X"fcb79ee3", X"00100793", X"70f601a3", X"10100737", X"70174783", X"01879793", X"4187d793",
        X"0607c263", X"01812403", X"01c12083", X"01412483", X"00200513", X"02010113", X"65c0006f", X"00000013",
        X"ea5ff06f", X"00000013", X"eb9ff06f", X"00000013", X"ecdff06f", X"00000013", X"eedff06f", X"00000013",
        X"f09ff06f", X"00000013", X"f25ff06f", X"00000013", X"f39ff06f", X"00000013", X"f4dff06f", X"00000013",
        X"f71ff06f", X"00000013", X"f8dff06f", X"ff010113", X"00812423", X"00050413", X"01855513", X"00112623",
        X"d7dff0ef", X"01045513", X"0ff57513", X"d71ff0ef", X"00845513", X"0ff57513", X"d65ff0ef", X"0ff47513",
        X"d5dff0ef", X"00812403", X"00c12083", X"02000513", X"01010113", X"5ec0006f", X"ff010113", X"00812423",
        X"00112623", X"00050413", X"00044503", X"00051a63", X"00c12083", X"00812403", X"01010113", X"00008067",
        X"00140413", X"5bc000ef", X"fe1ff06f", X"101007b7", X"10a79023", X"10b78123", X"101006b7", X"00a00793",
        X"1026c703", X"fff78793", X"fe079ce3", X"00008067", X"ff010113", X"00812423", X"00050413", X"00855513",
        X"00112623", X"00912223", X"00058493", X"cd1ff0ef", X"0ff47513", X"cc9ff0ef", X"00812403", X"00c12083",
        X"00048513", X"00412483", X"01010113", X"4940006f", X"f4010113", X"0a812c23", X"0b212823", X"0a112e23",
        X"0a912a23", X"0b312623", X"0b412423", X"0b512223", X"0b612023", X"09712e23", X"09812c23", X"09912a23",
        X"101007b7", X"00900713", X"10e78623", X"7d000413", X"10100937", X"10c94783", X"fff40413", X"fe041ce3",
        X"00200593", X"40000513", X"f45ff0ef", X"00000593", X"0000c537", X"f39ff0ef", X"00000593", X"00008537",
        X"f2dff0ef", X"00004537", X"00000593", X"05a50513", X"f1dff0ef", X"00000593", X"74200513", X"f11ff0ef",
        X"00200593", X"40000513", X"f05ff0ef", X"00100593", X"40000513", X"ef9ff0ef", X"00100593", X"40000513",
        X"eedff0ef", X"00100593", X"40000513", X"ee1ff0ef", X"00100593", X"40000513", X"ed5ff0ef", X"00c94783",
        X"01500713", X"0ff7f793", X"0037d793", X"00e79663", X"00100793", X"10f904a3", X"123457b7", X"67878793",
        X"10f02023", X"876547b7", X"32178793", X"10f02223", X"00100713", X"101007b7", X"10e781a3", X"00a00513",
        X"440000ef", X"00000a13", X"fff00c13", X"05500b13", X"101006b7", X"01010793", X"10068713", X"00300613",
        X"10002583", X"00478793", X"00b12623", X"1046a583", X"feb7ae23", X"00c70323", X"01870223", X"018702a3",
        X"09010593", X"fcb79ee3", X"00000993", X"01f00a93", X"02000b93", X"01010793", X"00f98533", X"fff00c93",
        X"fff00493", X"00000613", X"00000793", X"02fadc63", X"09849663", X"00198993", X"00400793", X"fcf99ce3",
        X"101007b7", X"00100713", X"10e783a3", X"001a0a13", X"f93a10e3", X"80001537", X"c9050513", X"2e4000ef",
        X"1480006f", X"00279713", X"00e50733", X"00074703", X"00178693", X"01670663", X"00068793", X"fb1ff06f",
        X"00078713", X"00070593", X"00170713", X"01770a63", X"00271693", X"00d506b3", X"0006c683", X"ff6684e3",
        X"40f586b3", X"00d65863", X"00058c93", X"00078493", X"00068613", X"00070793", X"f75ff06f", X"04600513",
        X"340000ef", X"0ff4f513", X"a95ff0ef", X"04c00513", X"330000ef", X"0ffcf513", X"a85ff0ef", X"02049a63",
        X"00900793", X"ff7c8913", X"0397cc63", X"409c87b3", X"00a00713", X"fff00913", X"02f75463", X"019484b3",
        X"01f4d913", X"00990933", X"40195913", X"0140006f", X"fd5c9ee3", X"01600793", X"00948913", X"fc97c8e3",
        X"04300513", X"2dc000ef", X"0ff97493", X"00048513", X"a2dff0ef", X"00a00513", X"2c8000ef", X"ef205ce3",
        X"101007b7", X"0ff9f993", X"10078793", X"00000713", X"00300613", X"fff00693", X"01378423", X"00c78323",
        X"00d78223", X"00d782a3", X"00170713", X"ff2748e3", X"04200513", X"28c000ef", X"0ffa7513", X"9e1ff0ef",
        X"04400513", X"27c000ef", X"00098513", X"9d1ff0ef", X"05000513", X"26c000ef", X"00048513", X"9c1ff0ef",
        X"00a00513", X"25c000ef", X"101007b7", X"00d00713", X"800024b7", X"10e78623", X"c0048493", X"0004a503",
        X"c0dff0ef", X"0004a783", X"80001537", X"ca450513", X"00178793", X"00f4a023", X"168000ef", X"0004a783",
        X"0017f793", X"10079a63", X"000054b7", X"5aa48493", X"00000793", X"000106b7", X"00179713", X"00f4c633",
        X"00e68733", X"00c71023", X"00178793", X"fed796e3", X"80001537", X"cac50513", X"128000ef", X"00000913",
        X"00010a37", X"01300b13", X"80001cb7", X"80001bb7", X"80001c37", X"00141793", X"00fa07b3", X"0084c9b3",
        X"0007da83", X"01099993", X"0109d993", X"03598a63", X"032b4663", X"01091513", X"cb4c8593", X"01055513",
        X"c11ff0ef", X"cb8b8593", X"00098513", X"c05ff0ef", X"c48c0593", X"000a8513", X"bf9ff0ef", X"00190913",
        X"00140413", X"fb4418e3", X"06090e63", X"80001537", X"cc050513", X"0ac000ef", X"00090513", X"b31ff0ef",
        X"00a00513", X"15c000ef", X"00042503", X"b21ff0ef", X"00442503", X"b19ff0ef", X"00842503", X"b11ff0ef",
        X"0b812403", X"0bc12083", X"0b412483", X"0b012903", X"0ac12983", X"0a812a03", X"0a412a83", X"0a012b03",
        X"09c12b83", X"09812c03", X"09412c83", X"00a00513", X"0c010113", X"10c0006f", X"000104b7", X"fff48493",
        X"ef1ff06f", X"0b812403", X"0bc12083", X"0b412483", X"0b012903", X"0ac12983", X"0a812a03", X"0a412a83",
        X"0a012b03", X"09c12b83", X"09812c03", X"09412c83", X"80001537", X"ccc50513", X"0c010113", X"0040006f",
        X"ff010113", X"00812423", X"00912223", X"00112623", X"00050493", X"00000413", X"008487b3", X"0007c503",
        X"00140413", X"00050663", X"098000ef", X"fedff06f", X"00d00513", X"08c000ef", X"00a00513", X"084000ef",
        X"00c12083", X"00040513", X"00812403", X"00412483", X"01010113", X"00008067", X"10000737", X"00c74783",
        X"01879693", X"00d74783", X"00e74503", X"00f74703", X"0ff7f793", X"01079793", X"0ff77713", X"00d7e7b3",
        X"0ff57513", X"00e7e7b3", X"00851513", X"00f56533", X"00008067", X"00000793", X"100006b7", X"fc800613",
        X"00a7c463", X"00008067", X"00c68323", X"0066c703", X"0ff77713", X"fe071ce3", X"00178793", X"fe5ff06f",
        X"800027b7", X"c047a783", X"ff010113", X"00812423", X"00112623", X"00050413", X"00078463", X"000780e7",
        X"10000737", X"01274783", X"0107f793", X"fe079ce3", X"0ff47413", X"00870823", X"00c12083", X"00812403",
        X"01010113", X"00008067", X"6c6c6548", X"6f77206f", X"2c646c72", X"34365520", X"2149492d", X"00000000",
        X"6967614d", X"000a2163", X"6c707061", X"74616369", X"0a6e6f69", X"00000000", X"6e6e7552", X"0a676e69",
        X"00000000", X"6b636f4c", X"0000000a", X"74706d45", X"77203b79", X"69746961", X"6620676e", X"4a20726f",
        X"20474154", X"67616d69", X"6f742065", X"6f6f6220", X"000a2e74", X"6967614d", X"00203a63", X"33323130",
        X"37363534", X"42413938", X"46454443", X"00000000", X"696c6143", X"74617262", X"206e6f69", X"6c696166",
        X"00006465", X"74697257", X"002e2e65", X"64616552", X"00002e2e", X"0000003a", X"203d2120", X"00000000",
        X"204d4152", X"6f727265", X"000a2e72", X"204d4152", X"21214b4f", X"0000000d", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000"

    );
end package;
