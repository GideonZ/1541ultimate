
library ieee;
use ieee.std_logic_1164.all;

package bootrom_pkg is
    type t_boot_data    is array(natural range <>) of std_logic_vector(31 downto 0);

    constant c_bootrom : t_boot_data(0 to 8191) := (
        X"30047073", X"01000117", X"ffc10113", X"00009197", X"03418193", X"00000517", X"16050513", X"30551073",
        X"34151073", X"30001073", X"30401073", X"34401073", X"32001073", X"30601073", X"b0001073", X"b8001073",
        X"b0201073", X"b8201073", X"00000093", X"00000213", X"00000293", X"00000313", X"00000393", X"00000813",
        X"00000893", X"00000913", X"00000993", X"00000a13", X"00000a93", X"00000b13", X"00000b93", X"00000c13",
        X"00000c93", X"00000d13", X"00000d93", X"00000e13", X"00000e93", X"00000f13", X"00000f93", X"00006597",
        X"7c058593", X"00008617", X"f5c60613", X"00008697", X"79468693", X"00d65c63", X"0005a703", X"00e62023",
        X"00458593", X"00460613", X"fedff06f", X"00008717", X"77470713", X"b0c18793", X"00f75863", X"00072023",
        X"00470713", X"ff5ff06f", X"00006997", X"d0898993", X"00006a17", X"d0ca0a13", X"0149da63", X"0009a303",
        X"000300e7", X"00498993", X"ff1ff06f", X"00000513", X"00000593", X"154000ef", X"34051073", X"00006997",
        X"ce098993", X"00006a17", X"cd8a0a13", X"0149da63", X"0009a303", X"000300e7", X"00498993", X"ff1ff06f",
        X"00000093", X"00008463", X"000080e7", X"10500073", X"0000006f", X"00000013", X"00000013", X"00000013",
        X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"ff810113", X"00812023", X"00912223",
        X"34202473", X"02044663", X"34102473", X"00041483", X"0034f493", X"00240413", X"34141073", X"00300413",
        X"00941863", X"34102473", X"00240413", X"34141073", X"10000437", X"04900493", X"00940fa3", X"00012403",
        X"00412483", X"00810113", X"30200073", X"ff010113", X"00812423", X"86018513", X"00112623", X"39d020ef",
        X"86018593", X"00812403", X"00c12083", X"00002537", X"82818613", X"77850513", X"01010113", X"0690406f",
        X"ff010113", X"00812423", X"88018513", X"00112623", X"2b9030ef", X"88018593", X"00812403", X"00c12083",
        X"00003537", X"82818613", X"28050513", X"01010113", X"0350406f", X"ff010113", X"00812423", X"89018513",
        X"00112623", X"5f9030ef", X"89018593", X"00812403", X"00c12083", X"00004537", X"82818613", X"fc450513",
        X"01010113", X"0010406f", X"ff010113", X"000097b7", X"00112623", X"8407a023", X"0d4000ef", X"00050613",
        X"000065b7", X"00006537", X"7d058593", X"7d850513", X"28d010ef", X"088000ef", X"00055c63", X"100007b7",
        X"02a00713", X"00e78823", X"00010537", X"7bc040ef", X"1c5040ef", X"00050593", X"02051663", X"00007537",
        X"010005b7", X"81850513", X"1dd040ef", X"00007537", X"000105b7", X"82450513", X"1cd040ef", X"00051a63",
        X"0000006f", X"00007537", X"83450513", X"231010ef", X"265040ef", X"00051c63", X"33d040ef", X"00055863",
        X"00007537", X"84c50513", X"261010ef", X"00c12083", X"00000513", X"01010113", X"00008067", X"10000737",
        X"00c74683", X"00d74783", X"00e74503", X"00f74703", X"01869693", X"01079793", X"00d7e7b3", X"00e7e7b3",
        X"00851513", X"00f56533", X"00008067", X"100007b7", X"00b7c503", X"00008067", X"10000737", X"02374783",
        X"02274503", X"02374683", X"00851513", X"00f56533", X"02274783", X"00879793", X"00d7e7b3", X"fef510e3",
        X"00008067", X"100007b7", X"ff000693", X"0127c703", X"01871713", X"41875713", X"00075863", X"0107c503",
        X"000788a3", X"00008067", X"fff50513", X"00a05a63", X"00d78323", X"0067c703", X"fe071ee3", X"fd1ff06f",
        X"ffe00513", X"00008067", X"000097b7", X"8407a783", X"ff010113", X"00812423", X"00112623", X"00050413",
        X"00078463", X"000780e7", X"10000737", X"01274783", X"0107f793", X"fe079ce3", X"0ff47413", X"00870823",
        X"00c12083", X"00812403", X"01010113", X"00008067", X"ff010113", X"00112623", X"5dc00513", X"f69ff0ef",
        X"fe055ce3", X"00c12083", X"01010113", X"00008067", X"ba010113", X"44812c23", X"44912a23", X"45212823",
        X"45312623", X"45412423", X"45512223", X"43712e23", X"43812c23", X"43912a23", X"43a12823", X"43b12623",
        X"44112e23", X"45612023", X"00050a13", X"00058a93", X"01900993", X"00000413", X"00100493", X"04300d93",
        X"00000913", X"00400b93", X"01800c13", X"00100c93", X"00200d13", X"01000b13", X"000d8663", X"000d8513",
        X"f29ff0ef", X"7d000513", X"eddff0ef", X"00054a63", X"07750863", X"04abc463", X"0b950a63", X"15a50e63",
        X"fffb0b13", X"fc0b1ae3", X"04300793", X"02fd8463", X"f41ff0ef", X"01800513", X"ef1ff0ef", X"01800513",
        X"ee9ff0ef", X"01800513", X"ee1ff0ef", X"ffe00413", X"03c0006f", X"01500d93", X"f9dff06f", X"fd8512e3",
        X"3e800513", X"e81ff0ef", X"fb851ce3", X"f05ff0ef", X"00600513", X"eb5ff0ef", X"fff00413", X"0100006f",
        X"ef1ff0ef", X"00600513", X"ea1ff0ef", X"45c12083", X"00040513", X"45812403", X"45412483", X"45012903",
        X"44c12983", X"44812a03", X"44412a83", X"44012b03", X"43c12b83", X"43812c03", X"43412c83", X"43012d03",
        X"42c12d83", X"46010113", X"00008067", X"08000b13", X"04300793", X"00fd9463", X"00100913", X"01810d93",
        X"012b0733", X"00a10c23", X"000d8693", X"00000793", X"00270713", X"3e800513", X"00e12623", X"00d12423",
        X"00f12223", X"de1ff0ef", X"06054c63", X"00812683", X"00412783", X"00c12703", X"00a680a3", X"00178793",
        X"00168693", X"fcf758e3", X"01a14783", X"01914703", X"fff7c793", X"0ff7f793", X"04f71463", X"04970863",
        X"fff48793", X"02f71e63", X"04090463", X"fff98993", X"0b304263", X"e1dff0ef", X"01800513", X"dcdff0ef",
        X"01800513", X"dc5ff0ef", X"01800513", X"dbdff0ef", X"ffd00413", X"f19ff06f", X"40000b13", X"f55ff06f",
        X"df1ff0ef", X"01500513", X"0700006f", X"02091c63", X"016d86b3", X"00000793", X"003dc603", X"001d8d93",
        X"00c787b3", X"0ff7f793", X"fedd98e3", X"410b0693", X"01010613", X"00c686b3", X"bfb6c683", X"fcf692e3",
        X"f89716e3", X"408a89b3", X"013b5463", X"000b0993", X"01305c63", X"008a0533", X"00098613", X"01b10593",
        X"0c0050ef", X"01340433", X"00148493", X"0ff4f493", X"01900993", X"00600513", X"d31ff0ef", X"00000d93",
        X"df5ff06f", X"fb010113", X"04812423", X"04912223", X"05212023", X"03512a23", X"03612823", X"03712623",
        X"03812423", X"03912223", X"04112623", X"03312e23", X"03412c23", X"03a12023", X"01b12e23", X"00050913",
        X"00058493", X"00c12623", X"00000413", X"00006ab7", X"00006b37", X"00006bb7", X"00006c37", X"05f00c93",
        X"04944063", X"04c12083", X"04812403", X"04412483", X"04012903", X"03c12983", X"03812a03", X"03412a83",
        X"03012b03", X"02c12b83", X"02812c03", X"02412c83", X"02012d03", X"01c12d83", X"05010113", X"00008067",
        X"00c12783", X"06078e63", X"00040593", X"dfcb0513", X"5cc010ef", X"00040d13", X"01040a13", X"069d5863",
        X"01a907b3", X"0007c583", X"e0cc0513", X"5b0010ef", X"001d0d13", X"ff4d14e3", X"40848d33", X"00000993",
        X"00890433", X"01000d93", X"03a98463", X"01340733", X"00074503", X"07f57513", X"fe050713", X"0ff77713",
        X"02ecec63", X"00198993", X"618010ef", X"fdb99ee3", X"00a00513", X"60c010ef", X"000a0413", X"f45ff06f",
        X"008905b3", X"e04a8513", X"f89ff06f", X"e14b8513", X"54c010ef", X"f9dff06f", X"02e00513", X"fc9ff06f",
        X"00100613", X"ec1ff06f", X"00154703", X"00054783", X"00871713", X"00f76733", X"00254783", X"00354503",
        X"01079793", X"00e7e7b3", X"01851513", X"00f56533", X"00008067", X"00050793", X"00c50633", X"0007c503",
        X"0005c703", X"00178793", X"00158593", X"40e50533", X"00c78463", X"fe0504e3", X"00008067", X"00c52783",
        X"ffe58593", X"ffe78793", X"02f5fa63", X"ff010113", X"00812423", X"00050413", X"00a55503", X"00112623",
        X"630040ef", X"02042783", X"00c12083", X"00812403", X"00f50533", X"01010113", X"00008067", X"00000513",
        X"00008067", X"00052703", X"00050693", X"02070463", X"00070793", X"02000513", X"03a00593", X"0007c603",
        X"00178793", X"02c57663", X"feb61ae3", X"00270613", X"00c78663", X"fff00513", X"00008067", X"00074603",
        X"03000713", X"fff00513", X"fee618e3", X"00f6a023", X"00000513", X"00008067", X"ff010113", X"00912223",
        X"00112623", X"00812423", X"00058493", X"02051263", X"00900513", X"00000793", X"00c12083", X"00812403",
        X"00f4a023", X"00412483", X"01010113", X"00008067", X"00052783", X"00050413", X"fc078ce3", X"0007c703",
        X"fc0708e3", X"00455683", X"0067d703", X"fce692e3", X"0017c503", X"681000ef", X"00157513", X"fa051ae3",
        X"00042783", X"fb5ff06f", X"02452783", X"04b78a63", X"ff010113", X"00812423", X"00912223", X"00112623",
        X"00050413", X"00058493", X"00058613", X"02850593", X"00154503", X"00100693", X"641000ef", X"00050663",
        X"00100513", X"fff00493", X"02942223", X"00c12083", X"00812403", X"00412483", X"01010113", X"00008067",
        X"00000513", X"00008067", X"ff010113", X"00812423", X"00912223", X"00112623", X"fff00793", X"000501a3",
        X"02f52223", X"00050493", X"f81ff0ef", X"00400413", X"06051c63", X"2274c783", X"2264c703", X"00300413",
        X"00879793", X"00e7e7b3", X"0000b737", X"a5570713", X"04e79c63", X"0284c783", X"0eb00713", X"00050413",
        X"00e78a63", X"01878793", X"0ff7f793", X"00100713", X"04f76863", X"000065b7", X"00300613", X"e1858593",
        X"05e48513", X"df1ff0ef", X"02050063", X"000065b7", X"00500613", X"e1c58593", X"07a48513", X"dd9ff0ef",
        X"00a03433", X"00141413", X"00c12083", X"00040513", X"00812403", X"00412483", X"01010113", X"00008067",
        X"00200413", X"fe5ff06f", X"fc010113", X"03212823", X"02112e23", X"02812c23", X"02912a23", X"03312623",
        X"03412423", X"03512223", X"03612023", X"01712e23", X"01812c23", X"01912a23", X"0005a023", X"00058913",
        X"de5ff0ef", X"2e054a63", X"000097b7", X"00251713", X"84478793", X"00e787b3", X"0007a403", X"00050493",
        X"00c00513", X"02040663", X"00892023", X"00044783", X"04079a63", X"0ff4f513", X"00040023", X"00a400a3",
        X"4a9000ef", X"00157793", X"00300513", X"04078863", X"03c12083", X"03812403", X"03412483", X"03012903",
        X"02c12983", X"02812a03", X"02412a83", X"02012b03", X"01c12b83", X"01812c03", X"01412c83", X"04010113",
        X"00008067", X"00144503", X"48d000ef", X"00157793", X"00000513", X"fa0790e3", X"fb9ff06f", X"00000593",
        X"00040513", X"e65ff0ef", X"00200713", X"00050793", X"06e51463", X"00010493", X"1ee40913", X"22e40a13",
        X"00048993", X"00090513", X"c81ff0ef", X"00a9a023", X"01090913", X"00498993", X"ff4916e3", X"01048913",
        X"00100993", X"0004a583", X"00300793", X"00058a63", X"00040513", X"e15ff0ef", X"00050793", X"02a9fc63",
        X"00448493", X"ff2490e3", X"00400713", X"00100513", X"00e79e63", X"f3dff06f", X"00400713", X"00100513",
        X"f2e788e3", X"00100713", X"00f77663", X"00d00513", X"f21ff06f", X"03444783", X"03344703", X"02442a03",
        X"00879793", X"00e7e7b3", X"20000713", X"fee790e3", X"03f44903", X"03e44783", X"00891913", X"00f96933",
        X"00091863", X"04c40513", X"be1ff0ef", X"00050913", X"03844983", X"01242823", X"00100713", X"fff98793",
        X"01340123", X"0ff7f793", X"faf762e3", X"03544c83", X"010c9793", X"0107d793", X"00f41523", X"f80788e3",
        X"fffc8793", X"0197f7b3", X"f80792e3", X"03a44b83", X"03944783", X"008b9b93", X"00fbebb3", X"01741423",
        X"00fbf793", X"f60794e3", X"03c44483", X"03b44783", X"00849493", X"00f4e4b3", X"00049863", X"04840513",
        X"b69ff0ef", X"00050493", X"03744a83", X"03644783", X"008a9a93", X"00faeab3", X"f20a8ae3", X"00090593",
        X"00098513", X"004bdc13", X"1e8040ef", X"015c0c33", X"00ac0c33", X"00050b13", X"f184eae3", X"418489b3",
        X"000c8593", X"00098513", X"1f4040ef", X"00050493", X"ef99eee3", X"100007b7", X"ff578793", X"eea7e8e3",
        X"000107b7", X"ff578793", X"0aa7fc63", X"00300993", X"00248493", X"015a0ab3", X"018a0c33", X"00942623",
        X"01442a23", X"01542c23", X"03842023", X"00300793", X"06f99063", X"05344783", X"05244703", X"00879793",
        X"00e7e7b3", X"00fbe7b3", X"ea0792e3", X"05440513", X"ab9ff0ef", X"00249793", X"1ff78793", X"00a42e23",
        X"0097d793", X"e8f964e3", X"80818713", X"00075783", X"01340023", X"00000513", X"00178793", X"01079793",
        X"0107d793", X"00f71023", X"00f41323", X"d85ff06f", X"e40b8ee3", X"00200713", X"015b0533", X"00149793",
        X"fae98ce3", X"009787b3", X"0017d793", X"0014f493", X"009787b3", X"fa5ff06f", X"00b00513", X"d55ff06f",
        X"000019b7", X"ff598993", X"00a9b9b3", X"00198993", X"f41ff06f", X"01b5c783", X"01a5c683", X"00050713",
        X"00879793", X"00d7e533", X"00300793", X"00f71e63", X"0155c783", X"0145c703", X"00879793", X"00e7e7b3",
        X"01079793", X"00f56533", X"00008067", X"00100793", X"14b7f063", X"00c52703", X"fe010113", X"00812c23",
        X"00912a23", X"00112e23", X"01212823", X"01312623", X"00050493", X"00058413", X"02e5fe63", X"00054703",
        X"00200693", X"0ad70463", X"00300693", X"0cd70a63", X"02f71263", X"0015d913", X"01852783", X"00b90933",
        X"00995593", X"00f585b3", X"b01ff0ef", X"02050463", X"fff00793", X"01c12083", X"01812403", X"01412483",
        X"01012903", X"00c12983", X"00078513", X"02010113", X"00008067", X"0184a783", X"00190993", X"0099d593",
        X"1ff97913", X"01248933", X"00f585b3", X"00048513", X"02894903", X"ab5ff0ef", X"fa051ce3", X"1ff9f993",
        X"013489b3", X"0289c783", X"00147413", X"00879793", X"0127e7b3", X"00040663", X"0047d793", X"f99ff06f",
        X"01479793", X"0147d793", X"f8dff06f", X"01852783", X"0085d593", X"00f585b3", X"a71ff0ef", X"f6051ae3",
        X"00141413", X"1fe47413", X"00848433", X"02944783", X"02844703", X"00879793", X"00e7e7b3", X"f59ff06f",
        X"01852783", X"0075d593", X"00f585b3", X"a3dff0ef", X"f40510e3", X"00241413", X"02848513", X"1fc47413",
        X"00850533", X"8c5ff0ef", X"00451793", X"f8dff06f", X"00100793", X"00078513", X"00008067", X"fd010113",
        X"00852583", X"02812423", X"02912223", X"02112623", X"03212023", X"01312e23", X"00052823", X"00052403",
        X"00050493", X"06059063", X"00044703", X"00200793", X"00e7f663", X"01c42783", X"04079863", X"00845783",
        X"02079263", X"00200513", X"02c12083", X"02812403", X"02412483", X"02012903", X"01c12983", X"03010113",
        X"00008067", X"01c42503", X"00a4ac23", X"00b4aa23", X"fc050ae3", X"02840413", X"0084ae23", X"00000513",
        X"fc9ff06f", X"00058793", X"00a45703", X"00078593", X"fff00913", X"00100993", X"02071263", X"0004a503",
        X"e0dff0ef", X"00050593", X"03250463", X"f8a9fce3", X"00c42783", X"fef564e3", X"f8dff06f", X"00040513",
        X"00f12623", X"839ff0ef", X"00c12583", X"f9dff06f", X"00100513", X"f75ff06f", X"fe010113", X"01212823",
        X"01052903", X"00812c23", X"00912a23", X"00112e23", X"01312623", X"02090913", X"002007b7", X"00052483",
        X"00050413", X"00f96463", X"00052c23", X"01842783", X"00400513", X"02078863", X"1ff97993", X"08099a63",
        X"01442583", X"00178793", X"00f42c23", X"02059a63", X"0084d703", X"00595793", X"06e7ec63", X"00042c23",
        X"00400513", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"02010113", X"00008067",
        X"00a4d783", X"00995713", X"fff78793", X"00e7f7b3", X"04079063", X"00048513", X"d35ff0ef", X"00050593",
        X"00100793", X"00200513", X"fab7fee3", X"fff00793", X"00100513", X"faf588e3", X"00c4a783", X"faf5f0e3",
        X"00b42a23", X"00048513", X"f54ff0ef", X"00a42c23", X"02848493", X"013484b3", X"01242823", X"00942e23",
        X"00000513", X"f81ff06f", X"fd010113", X"01512a23", X"00052a83", X"02912223", X"03212023", X"02112623",
        X"02812423", X"01312e23", X"01412c23", X"01612823", X"01712623", X"01812423", X"00050493", X"00058913",
        X"02f00693", X"05c00713", X"00094783", X"08d78263", X"08e78063", X"0004a423", X"00094703", X"01f00793",
        X"06e7fc63", X"00006a37", X"02048993", X"00006b37", X"e34a0a13", X"028a8b93", X"00b00613", X"02000593",
        X"00098513", X"6e4040ef", X"00000693", X"00000713", X"00800613", X"02000813", X"02f00893", X"05c00313",
        X"02e00e13", X"00b00e93", X"01900f13", X"00170713", X"00e907b3", X"fff7c783", X"06f87863", X"01178463",
        X"0e679c63", X"02f00513", X"05c00593", X"04c0006f", X"00190913", X"f75ff06f", X"02812403", X"f8000793",
        X"02c12083", X"02012903", X"01c12983", X"01812a03", X"01412a83", X"01012b03", X"00c12b83", X"00812c03",
        X"02f485a3", X"00048513", X"02412483", X"03010113", X"d2dff06f", X"00170713", X"00e90633", X"00064603",
        X"fea60ae3", X"feb608e3", X"00e90933", X"0a068e63", X"0204c683", X"0e500713", X"00e69663", X"00500713",
        X"02e48023", X"0217b793", X"00279793", X"02f485a3", X"00048513", X"0004ac03", X"ce5ff0ef", X"00050413",
        X"08051e63", X"0184a583", X"000c0513", X"edcff0ef", X"00050413", X"08051463", X"01c4a503", X"00054783",
        X"06078c63", X"00b54783", X"03f7f793", X"00f48323", X"00b54783", X"0087f793", X"00079a63", X"00b00613",
        X"00098593", X"d70ff0ef", X"04050a63", X"00048513", X"d69ff0ef", X"fa9ff06f", X"0dc78463", X"02c6f663",
        X"01879593", X"4185d593", X"0005d863", X"07f7f793", X"00fa07b3", X"0007c783", X"e24b0593", X"0005c503",
        X"0a050863", X"00a79663", X"00600413", X"0280006f", X"00158593", X"fe9ff06f", X"00400413", X"02b4c783",
        X"04040463", X"00400713", X"00e41663", X"0047f793", X"06078463", X"02c12083", X"00040513", X"02812403",
        X"02412483", X"02012903", X"01c12983", X"01812a03", X"01412a83", X"01012b03", X"00c12b83", X"00812c03",
        X"03010113", X"00008067", X"0047f793", X"fc0794e3", X"0064c783", X"0107f793", X"02078063", X"0104a583",
        X"000ac503", X"1ff5f593", X"00bb85b3", X"a49ff0ef", X"00a4a423", X"e05ff06f", X"00500413", X"f99ff06f",
        X"f7d604e3", X"00800693", X"00b00613", X"e21ff06f", X"f9f78593", X"0ff5f593", X"00bf6663", X"fe078793",
        X"0ff7f793", X"00d985b3", X"00f58023", X"00168693", X"dfdff06f", X"fd010113", X"00a12623", X"01c10513",
        X"02812423", X"02112623", X"00b12423", X"00060413", X"00b12e23", X"cb0ff0ef", X"04054e63", X"000097b7",
        X"84478713", X"00251513", X"00a70733", X"00072703", X"84478793", X"00070463", X"00070023", X"00c12703",
        X"00070463", X"00070023", X"00a787b3", X"00e7a023", X"00000513", X"00040863", X"00c10593", X"00810513",
        X"e48ff0ef", X"02c12083", X"02812403", X"03010113", X"00008067", X"00b00513", X"fedff06f", X"fa010113",
        X"04912a23", X"04112e23", X"04812c23", X"05212823", X"05312623", X"05412423", X"00b12623", X"00900493",
        X"08050863", X"00050413", X"01010593", X"00c10513", X"00060913", X"df4ff0ef", X"00050493", X"08051e63",
        X"01012983", X"00c12583", X"01410513", X"01312a23", X"c79ff0ef", X"00050493", X"08051063", X"03f10783",
        X"0607ca63", X"01a14783", X"0107f793", X"06079a63", X"03012a03", X"0009c503", X"00197913", X"000a0593",
        X"8f5ff0ef", X"00a42423", X"01ca0513", X"b1cff0ef", X"0069d783", X"00a42623", X"01342023", X"00f41223",
        X"01240823", X"000408a3", X"00042e23", X"00042a23", X"05c12083", X"05812403", X"05012903", X"04c12983",
        X"04812a03", X"00048513", X"05412483", X"06010113", X"00008067", X"00600493", X"00042023", X"fd5ff06f",
        X"00400493", X"ff5ff06f", X"fb010113", X"04812423", X"04912223", X"05212023", X"03312e23", X"03412c23",
        X"04112623", X"03512a23", X"03612823", X"03712623", X"03812423", X"03912223", X"03a12023", X"00058993",
        X"0006a023", X"01c10593", X"00050493", X"00060913", X"00068a13", X"b64ff0ef", X"00050413", X"08051463",
        X"0114c783", X"00078413", X"06079e63", X"0104c783", X"00700413", X"0017f793", X"06078663", X"00c4a403",
        X"0144a783", X"40f40433", X"00897463", X"00090413", X"20000b13", X"02048a93", X"1ff00b93", X"fff00c13",
        X"04040263", X"0144a783", X"1ff7f713", X"12071663", X"01c12d03", X"0097d713", X"00ad5c83", X"fffc8c93",
        X"00ecfcb3", X"080c9263", X"04079c63", X"0084a503", X"00100793", X"04a7ee63", X"00200793", X"00f488a3",
        X"00200413", X"04c12083", X"00040513", X"04812403", X"04412483", X"04012903", X"03c12983", X"03812a03",
        X"03412a83", X"03012b03", X"02c12b83", X"02812c03", X"02412c83", X"02012d03", X"05010113", X"00008067",
        X"0184a583", X"0004a503", X"fa4ff0ef", X"fa5ff06f", X"01851a63", X"00100793", X"00f488a3", X"00100413",
        X"fa5ff06f", X"00a4ac23", X"0184a583", X"000d0513", X"9ccff0ef", X"f80502e3", X"00ac8633", X"048bfa63",
        X"00ad5783", X"00945913", X"012c8733", X"00e7f463", X"41978933", X"001d4503", X"00090693", X"00098593",
        X"118000ef", X"fa0518e3", X"00991793", X"000a2703", X"40f40433", X"00f989b3", X"00f70733", X"00ea2023",
        X"0144a703", X"00f707b3", X"00f4aa23", X"ef5ff06f", X"01c4a783", X"02c78063", X"001d4503", X"00100693",
        X"000a8593", X"00c12623", X"0d0000ef", X"00c12603", X"f60512e3", X"00c4ae23", X"0144a683", X"1ff6f693",
        X"40db07b3", X"00f47463", X"00040793", X"00000713", X"00e68633", X"00ca8633", X"00064583", X"00e98633",
        X"00170713", X"00b60023", X"fee794e3", X"f81ff06f", X"fe010113", X"00c10593", X"00812c23", X"00112e23",
        X"00050413", X"994ff0ef", X"00051463", X"00042023", X"01c12083", X"01812403", X"02010113", X"00008067",
        X"02051063", X"8101c683", X"00069863", X"00100693", X"8001ac23", X"80d18823", X"8181a503", X"00008067",
        X"00000513", X"00008067", X"ff010113", X"00112623", X"fd1ff0ef", X"00050863", X"00c12083", X"01010113",
        X"45d0006f", X"00c12083", X"00300513", X"01010113", X"00008067", X"fd5ff06f", X"fe010113", X"00112e23",
        X"00b12623", X"00c12423", X"00d12223", X"f95ff0ef", X"00050e63", X"00412683", X"00812603", X"00c12583",
        X"01c12083", X"02010113", X"4310006f", X"01c12083", X"00300513", X"02010113", X"00008067", X"000097b7",
        X"01000737", X"83078793", X"b0c18693", X"00070713", X"00050613", X"0007a503", X"02e68063", X"00c506b3",
        X"00e6f863", X"00c686b3", X"00d7a023", X"00008067", X"00e7a023", X"00008067", X"00000513", X"00008067",
        X"ff010113", X"00812423", X"00112623", X"00a00793", X"00050413", X"00f51663", X"00d00513", X"b6dfe0ef",
        X"00040513", X"00812403", X"00c12083", X"01010113", X"b59fe06f", X"00006737", X"00c58633", X"f1870713",
        X"00f57793", X"00f707b3", X"0007c783", X"fff60613", X"40455513", X"00f60023", X"fec594e3", X"00008067",
        X"ee010113", X"11612023", X"00006b37", X"0f712e23", X"0f812c23", X"ebcb0793", X"00006bb7", X"00006c37",
        X"10812c23", X"11212823", X"11312623", X"11412423", X"0fa12823", X"10112e23", X"10912a23", X"11512223",
        X"0f912a23", X"0fb12623", X"00050993", X"00058a13", X"00060913", X"00068413", X"00000d13", X"00f12223",
        X"eb4b8b93", X"f18c0c13", X"00094503", X"04051263", X"11c12083", X"11812403", X"11412483", X"11012903",
        X"10c12983", X"10812a03", X"10412a83", X"10012b03", X"0fc12b83", X"0f812c03", X"0f412c83", X"0ec12d83",
        X"000d0513", X"0f012d03", X"12010113", X"00008067", X"02500793", X"3af51a63", X"00194c83", X"03000713",
        X"00290793", X"08ec8e63", X"02d00713", X"00ec9663", X"00294c83", X"00390793", X"02300713", X"00178913",
        X"08ec9a63", X"0007cc83", X"00042483", X"00000693", X"00440413", X"07800793", X"0197ee63", X"06100793",
        X"0797ee63", X"04200793", X"28fc8c63", X"05800793", X"24fc8263", X"000a0593", X"02500513", X"000980e7",
        X"000a0593", X"000c8513", X"000980e7", X"002d0d13", X"f39ff06f", X"00249793", X"009787b3", X"fff64c83",
        X"00179793", X"00f704b3", X"00060913", X"fd0c8713", X"0ff77793", X"00190613", X"fcf5fee3", X"f99ff06f",
        X"00100693", X"00078913", X"00000493", X"00900593", X"fddff06f", X"00000693", X"fedff06f", X"f9ec8793",
        X"0ff7f793", X"01600713", X"f8f766e3", X"00412703", X"00279793", X"00e787b3", X"0007a783", X"00078067",
        X"07500713", X"00042783", X"00440a93", X"01010d93", X"06ec8863", X"0607d663", X"02d00713", X"06e10023",
        X"40f007b3", X"06110b13", X"00100413", X"000d8c93", X"00a00593", X"00078513", X"00d12623", X"00f12423",
        X"484030ef", X"00ac0533", X"00054603", X"00812783", X"00a00593", X"00cc8023", X"00078513", X"420030ef",
        X"00812603", X"00900813", X"001c8c93", X"00c12683", X"00140413", X"00050793", X"fac86ce3", X"0280006f",
        X"00078863", X"06010b13", X"00000413", X"fa1ff06f", X"03000793", X"00f10823", X"06010b13", X"00100413",
        X"01110c93", X"04068263", X"408486b3", X"00000613", X"0084c463", X"00068613", X"000c8513", X"03000593",
        X"00c12423", X"00d12623", X"561030ef", X"00812603", X"00000793", X"00cc8cb3", X"0084c663", X"00c12683",
        X"00068793", X"00f40433", X"000b0693", X"000c8793", X"0140006f", X"fff7c603", X"fff78793", X"00168693",
        X"fec68fa3", X"ffb798e3", X"40fc8cb3", X"019b0733", X"00070023", X"0a945e63", X"408484b3", X"00000d93",
        X"06010c93", X"0480006f", X"00042c83", X"00440a93", X"000c9463", X"000b8c93", X"00000413", X"0080006f",
        X"00140413", X"008c87b3", X"0007c783", X"fe079ae3", X"40848db3", X"00944663", X"00000d93", X"00048863",
        X"0084d463", X"00048413", X"00000493", X"00048793", X"0e00006f", X"00044503", X"00440493", X"000a0593",
        X"000980e7", X"001d0d13", X"00048413", X"d3dff06f", X"00042503", X"00800613", X"06010593", X"00440a93",
        X"c95ff0ef", X"00000d93", X"00000493", X"00800413", X"f71ff06f", X"00440a93", X"0c048e63", X"00042503",
        X"00048613", X"06010593", X"c6dff0ef", X"00048413", X"00000d93", X"00000493", X"f49ff06f", X"00042503",
        X"00200613", X"06010593", X"00440a93", X"c49ff0ef", X"00000d93", X"00000493", X"00200413", X"f25ff06f",
        X"00042783", X"00440a93", X"00800493", X"0017f713", X"fff48493", X"02a00693", X"00071463", X"02e00693",
        X"06010713", X"00970733", X"00d70023", X"4017d793", X"fc049ee3", X"00000d93", X"f75ff06f", X"000a0593",
        X"02000513", X"00f12423", X"000980e7", X"00812783", X"fff00713", X"fff78793", X"fee792e3", X"009d04b3",
        X"008c8d33", X"419d07b3", X"02f04c63", X"00045463", X"00000413", X"00940433", X"000d8493", X"02904c63",
        X"000dd463", X"00000d93", X"008d8d33", X"000a8413", X"c39ff06f", X"00000d93", X"00000413", X"e85ff06f",
        X"000cc503", X"000a0593", X"001c8c93", X"000980e7", X"fb5ff06f", X"000a0593", X"02000513", X"000980e7",
        X"fff48493", X"fb9ff06f", X"000a0593", X"00190913", X"000980e7", X"001d0d13", X"bf1ff06f", X"fc010113",
        X"02c12423", X"00050613", X"00002537", X"02b12223", X"02d12623", X"00000593", X"02410693", X"84050513",
        X"00112e23", X"02e12823", X"02f12a23", X"03012c23", X"03112e23", X"00d12623", X"b49ff0ef", X"01c12083",
        X"04010113", X"00008067", X"ff010113", X"00812423", X"00912223", X"00112623", X"00050493", X"00000413",
        X"008487b3", X"0007c503", X"00140413", X"02051663", X"00d00513", X"e34fe0ef", X"00a00513", X"e2cfe0ef",
        X"00c12083", X"00040513", X"00812403", X"00412483", X"01010113", X"00008067", X"e10fe0ef", X"fc5ff06f",
        X"ff010113", X"00812423", X"00000593", X"00050413", X"0ff57513", X"00112623", X"a69ff0ef", X"00c12083",
        X"00040513", X"00812403", X"01010113", X"00008067", X"00008067", X"00052783", X"00c7a783", X"00078067",
        X"00200513", X"00008067", X"00300513", X"00008067", X"00300513", X"00008067", X"00800593", X"43d0206f",
        X"000067b7", X"f3478793", X"00f52023", X"00052223", X"00008067", X"ff010113", X"00812423", X"00050413",
        X"00042a23", X"00042823", X"00b42423", X"00c42023", X"00042223", X"00060513", X"00112623", X"401020ef",
        X"00c12083", X"00a42623", X"00812403", X"01010113", X"00008067", X"fc010113", X"02912a23", X"00050493",
        X"00052503", X"03212823", X"03412423", X"02112e23", X"00058a13", X"02812c23", X"03312623", X"03512223",
        X"03612023", X"01712e23", X"01812c23", X"01912a23", X"01a12823", X"3a9020ef", X"00050913", X"0084a503",
        X"00100693", X"000a0613", X"00052783", X"00090593", X"0107a783", X"000780e7", X"04050463", X"00090513",
        X"381020ef", X"ffe00513", X"03c12083", X"03812403", X"03412483", X"03012903", X"02c12983", X"02812a03",
        X"02412a83", X"02012b03", X"01c12b83", X"01812c03", X"01412c83", X"01012d03", X"04010113", X"00008067",
        X"1ff94783", X"1fe94703", X"00879793", X"00e7e7b3", X"0000b737", X"a5570713", X"00e78a63", X"00090513",
        X"321020ef", X"ffd00513", X"fa1ff06f", X"1be90413", X"04200593", X"00040513", X"889fe0ef", X"1fe90a93",
        X"00006b37", X"00f00b93", X"00500c13", X"00444683", X"08068063", X"00944703", X"00844783", X"00b44983",
        X"00871713", X"00f76733", X"00a44783", X"01899993", X"00f44c83", X"01079793", X"00e7e7b3", X"00d44703",
        X"00f9e9b3", X"00c44783", X"00871713", X"018c9c93", X"00f76733", X"00e44783", X"00098593", X"f50b0513",
        X"01079793", X"00e7e7b3", X"00fcecb3", X"000c8613", X"d4dff0ef", X"00444703", X"013a09b3", X"01770463",
        X"03871663", X"00098593", X"00048513", X"e89ff0ef", X"01040413", X"f68a9ce3", X"00090513", X"00100593",
        X"259020ef", X"00000513", X"ee1ff06f", X"01400513", X"00e12623", X"241020ef", X"00c12703", X"0084a583",
        X"000c8693", X"00098613", X"00050d13", X"398000ef", X"0104a783", X"00078e63", X"01a7a823", X"0044a783",
        X"01a4a823", X"00178793", X"00f4a223", X"fa5ff06f", X"01a4aa23", X"fe9ff06f", X"fb010113", X"04812423",
        X"00050413", X"00852503", X"04912223", X"04112623", X"00052783", X"05212023", X"03312e23", X"0087a783",
        X"03412c23", X"03512a23", X"03612823", X"03712623", X"03812423", X"03912223", X"00058493", X"000780e7",
        X"fff00793", X"04051663", X"00842503", X"00c42583", X"00100693", X"00052783", X"00000613", X"0107a783",
        X"000780e7", X"ffe00793", X"02051463", X"08048463", X"00842503", X"01c10613", X"00100593", X"00052783",
        X"0187a783", X"000780e7", X"04050063", X"ffd00793", X"04c12083", X"04812403", X"04412483", X"04012903",
        X"03c12983", X"03812a03", X"03412a83", X"03012b03", X"02c12b83", X"02812c03", X"02412c83", X"00078513",
        X"05010113", X"00008067", X"01400513", X"129020ef", X"00050493", X"00100713", X"01c12683", X"00842583",
        X"00000613", X"280000ef", X"00942a23", X"00100793", X"fa1ff06f", X"00c42783", X"1ff7c703", X"1fe7c683",
        X"00871713", X"00d76733", X"0000b6b7", X"a5568693", X"02d70a63", X"00842503", X"01c10613", X"00100593",
        X"00052783", X"0187a783", X"000780e7", X"f60510e3", X"01400513", X"0c1020ef", X"00050493", X"00000713",
        X"f99ff06f", X"0377c703", X"0367c683", X"010005b7", X"00871713", X"00d76733", X"0387c683", X"fff58593",
        X"00544637", X"01069693", X"00e6e6b3", X"0397c703", X"14660613", X"01871713", X"00d76733", X"00b77733",
        X"04c71e63", X"00842503", X"01c10613", X"00100593", X"00052783", X"0187a783", X"000780e7", X"00050663",
        X"ffc00793", X"eedff06f", X"01400513", X"049020ef", X"01c12683", X"00842583", X"00600713", X"00000613",
        X"00050493", X"1a0000ef", X"00006537", X"00942a23", X"f7450513", X"b35ff0ef", X"f15ff06f", X"0537c683",
        X"0527c703", X"00869693", X"00e6e6b3", X"0547c703", X"0557c783", X"01071713", X"00d76733", X"01879793",
        X"00e7e7b3", X"00b7f7b3", X"02c79a63", X"00842503", X"01c10613", X"00100593", X"00052783", X"0187a783",
        X"000780e7", X"f6051ee3", X"01400513", X"7c8020ef", X"00050493", X"00c00713", X"ea1ff06f", X"01442583",
        X"00006537", X"f8c50513", X"a75ff0ef", X"00c42a03", X"00042223", X"00006ab7", X"1bea0493", X"00f00b13",
        X"1fea0a13", X"00006bb7", X"00500c13", X"00006cb7", X"0044c683", X"08068463", X"0094c703", X"0084c783",
        X"00b4c903", X"00871713", X"00f76733", X"00a4c783", X"01891913", X"00f4c603", X"01079793", X"00e7e7b3",
        X"00d4c703", X"00f96933", X"00c4c783", X"00871713", X"01861613", X"00f76733", X"00e4c783", X"00090593",
        X"fc4a8513", X"01079793", X"00e7e7b3", X"00f66633", X"00c12e23", X"9e9ff0ef", X"0044c703", X"01670463",
        X"03871663", X"00090593", X"00040513", X"b29ff0ef", X"00050593", X"fe8b8513", X"9c5ff0ef", X"01048493",
        X"f69a18e3", X"00442783", X"d89ff06f", X"01400513", X"00e12623", X"6e0020ef", X"00c12703", X"01c12683",
        X"00842583", X"00090613", X"00050993", X"038000ef", X"00098593", X"004c8513", X"985ff0ef", X"01042783",
        X"00078e63", X"0137a823", X"00442783", X"01342823", X"00178793", X"00f42223", X"fa5ff06f", X"01342a23",
        X"fe9ff06f", X"00050793", X"0007a823", X"00b7a023", X"00c7a223", X"00d7a423", X"00e78623", X"00058513",
        X"00069c63", X"0005a703", X"00878613", X"00100593", X"01872703", X"00070067", X"00008067", X"00052503",
        X"00050863", X"00052783", X"00c7a783", X"00078067", X"00100513", X"00008067", X"00050793", X"00052503",
        X"02050063", X"0087a703", X"02e67063", X"0047a703", X"00052783", X"00e60633", X"0107a783", X"00078067",
        X"00300513", X"00008067", X"00400513", X"00008067", X"00100713", X"00e59a63", X"00852703", X"00000513",
        X"00e62023", X"00008067", X"00052503", X"00050863", X"00052783", X"0187a783", X"00078067", X"00300513",
        X"00008067", X"00008067", X"00000513", X"00008067", X"00006537", X"01c50513", X"00008067", X"00008067",
        X"00000513", X"00008067", X"00008067", X"00008067", X"00008067", X"00100513", X"00008067", X"20000513",
        X"00008067", X"00100513", X"00008067", X"00000513", X"00008067", X"fff00513", X"00008067", X"00000513",
        X"00008067", X"00052783", X"0387a783", X"00078067", X"00000513", X"00008067", X"00000513", X"00008067",
        X"20000513", X"00008067", X"00000513", X"00008067", X"00068513", X"00065463", X"00000613", X"0ff00593",
        X"3480306f", X"00008067", X"00008067", X"00008067", X"00000513", X"00008067", X"00008067", X"00008067",
        X"00008067", X"ff010113", X"00812423", X"00050413", X"00052503", X"00112623", X"00050463", X"504020ef",
        X"00842503", X"00050a63", X"00812403", X"00c12083", X"01010113", X"4ec0206f", X"00c12083", X"00812403",
        X"01010113", X"00008067", X"00400593", X"4cc0206f", X"ff010113", X"00912223", X"00812423", X"01000513",
        X"84c18413", X"00112623", X"00042223", X"4b0020ef", X"00a42023", X"00400513", X"4a4020ef", X"00400793",
        X"00a42423", X"00f42623", X"00042823", X"00812403", X"00c12083", X"00100713", X"84c18593", X"00412483",
        X"82e18023", X"00002537", X"82818613", X"54450513", X"01010113", X"4700206f", X"fe010113", X"01312623",
        X"8201c783", X"00112e23", X"00812c23", X"00912a23", X"01212823", X"01412423", X"00079463", X"f75ff0ef",
        X"00000913", X"84c18413", X"01042783", X"0ef94263", X"00400513", X"420020ef", X"000067b7", X"02c78793",
        X"00f52023", X"8201c783", X"00050493", X"00079463", X"f41ff0ef", X"01042a03", X"00c42783", X"06fa1263",
        X"01000913", X"000a0463", X"001a1913", X"01242623", X"200007b7", X"fff00513", X"00f97463", X"00291513",
        X"3dc020ef", X"00050993", X"00090513", X"3d0020ef", X"00050913", X"00842683", X"00042503", X"00000793",
        X"0947ce63", X"00050463", X"3b8020ef", X"00842503", X"00050463", X"3ac020ef", X"01342023", X"01242423",
        X"01042703", X"00042783", X"00271693", X"00d787b3", X"0097a023", X"00842783", X"00e787b3", X"00078023",
        X"01042783", X"00178793", X"00f42823", X"01c12083", X"01812403", X"01012903", X"00c12983", X"00812a03",
        X"00048513", X"01412483", X"02010113", X"00008067", X"00042783", X"00291713", X"00e787b3", X"0007a483",
        X"0004a783", X"00048513", X"0087a783", X"000780e7", X"fa051ee3", X"00190913", X"ef1ff06f", X"00279713",
        X"00e50633", X"00062603", X"00e98733", X"00c72023", X"00f68733", X"00074603", X"00f90733", X"00178793",
        X"00c70023", X"f3dff06f", X"01052503", X"00008067", X"00000513", X"00008067", X"00008067", X"ff010113",
        X"000067b7", X"00058713", X"00112623", X"00060513", X"12c78593", X"0ff00693", X"0005c783", X"00d79c63",
        X"01000613", X"79d020ef", X"00c12083", X"01010113", X"00008067", X"fee786e3", X"01058593", X"fddff06f",
        X"100607b7", X"00100713", X"20e78423", X"00300713", X"20e78023", X"4105d713", X"0ff77713", X"20e78023",
        X"4085d713", X"0ff77713", X"20e78023", X"0ff5f593", X"20b78023", X"10060737", X"00000793", X"00c7ca63",
        X"100607b7", X"00300713", X"20e78423", X"00008067", X"20074503", X"00f685b3", X"00178793", X"00a58023",
        X"fddff06f", X"00452503", X"00008067", X"00852583", X"00452503", X"ff010113", X"00112623", X"654020ef",
        X"00c12083", X"01010113", X"00008067", X"ff010113", X"000067b7", X"00112623", X"00812423", X"12c78793",
        X"0ff00813", X"0007c703", X"01071663", X"00000413", X"02c0006f", X"02b71e63", X"00c7a403", X"0086d463",
        X"00068413", X"00052703", X"0087a583", X"00060693", X"01c72703", X"00040613", X"000700e7", X"00c12083",
        X"00040513", X"00812403", X"01010113", X"00008067", X"01078793", X"fb1ff06f", X"fe010113", X"00912a23",
        X"00058493", X"00452583", X"00812c23", X"00050413", X"00048513", X"00112e23", X"01212823", X"00c12623",
        X"00d12423", X"00b12223", X"5cc020ef", X"01442783", X"00412583", X"00f51933", X"00048513", X"63c020ef",
        X"00042783", X"00a965b3", X"00040513", X"01812403", X"00812683", X"00c12603", X"01c12083", X"01412483",
        X"01012903", X"01c7a783", X"02010113", X"00078067", X"100607b7", X"00100713", X"20e78423", X"07700713",
        X"20e78023", X"20078023", X"20078023", X"20078023", X"04000713", X"20078793", X"fff00693", X"00d78023",
        X"fff70713", X"fe071ce3", X"00000793", X"10060737", X"04000693", X"20074503", X"00f58633", X"00178793",
        X"00a60023", X"fed798e3", X"00300793", X"20f70423", X"00008067", X"00052783", X"0287a783", X"00078067",
        X"01000513", X"00008067", X"01852703", X"00052783", X"00e585b3", X"01452703", X"01c7a783", X"00e595b3",
        X"00078067", X"00052783", X"01852703", X"0407a783", X"00e585b3", X"00078067", X"01452783", X"00100693",
        X"00452703", X"00f595b3", X"100607b7", X"20d78423", X"00300693", X"20d78023", X"4105d693", X"0ff6f693",
        X"20d78023", X"4085d693", X"0ff6f693", X"20d78023", X"0ff5f593", X"20b78023", X"40275713", X"00000793",
        X"100605b7", X"00e7cc63", X"100607b7", X"00300713", X"20e78423", X"00100513", X"00008067", X"2005a503",
        X"00279693", X"00d606b3", X"00a6a023", X"00178793", X"fd5ff06f", X"01452783", X"00100713", X"00f595b3",
        X"100607b7", X"20e78423", X"00300713", X"20e78023", X"4105d713", X"0ff77713", X"20e78023", X"4085d713",
        X"0ff77713", X"20e78023", X"0ff5f593", X"20b78023", X"20060713", X"2007a683", X"00460613", X"fed62e23",
        X"fec71ae3", X"00300713", X"20e78423", X"00100513", X"00008067", X"00058793", X"00852583", X"ff010113",
        X"00078513", X"00112623", X"3ec020ef", X"00c12083", X"01010113", X"00008067", X"100607b7", X"00100713",
        X"20e78423", X"3d2a8737", X"f9a70713", X"20e7a023", X"00300713", X"20e78423", X"00008067", X"100607b7",
        X"00100713", X"20e78423", X"3d2a8737", X"fa970713", X"20e7a023", X"00300713", X"20e78423", X"00008067",
        X"02000593", X"7350106f", X"fc010113", X"02912a23", X"00058493", X"00452583", X"02812c23", X"00050413",
        X"00048513", X"02112e23", X"03212823", X"00b12623", X"364020ef", X"01442783", X"00c12583", X"00006937",
        X"00f51433", X"00048513", X"3d0020ef", X"000065b7", X"00a46433", X"01400613", X"11858593", X"01c10513",
        X"3c1020ef", X"01041713", X"01075713", X"00841793", X"00875713", X"00e7e7b3", X"41045413", X"02f11023",
        X"00300793", X"028102a3", X"02f10223", X"00000413", X"01400493", X"01c10793", X"008787b3", X"0007c583",
        X"09c90513", X"00140413", X"954ff0ef", X"fe9414e3", X"100607b7", X"60078223", X"60078223", X"10060737",
        X"00000793", X"01400693", X"01c10613", X"00f60633", X"00064603", X"00178793", X"60c70423", X"fed796e3",
        X"60070223", X"60070223", X"03c12083", X"03812403", X"03412483", X"03012903", X"04010113", X"00008067",
        X"fe010113", X"00812c23", X"00050413", X"00c52503", X"00112e23", X"00912a23", X"625010ef", X"10060737",
        X"00100793", X"20f70423", X"323237b7", X"23278793", X"20f72023", X"00c42703", X"00000793", X"100606b7",
        X"06e7ca63", X"100604b7", X"00300793", X"20f48423", X"00c42583", X"00a12623", X"b69fd0ef", X"00100793",
        X"20f48423", X"00c42703", X"353537b7", X"00c12503", X"53578793", X"20f4a023", X"100606b7", X"00000793",
        X"04e7c463", X"100607b7", X"00300713", X"20e78423", X"00c42583", X"00a12623", X"b29fd0ef", X"01812403",
        X"00c12503", X"01c12083", X"01412483", X"02010113", X"5910106f", X"2006c583", X"00f50633", X"00178793",
        X"00b60023", X"f7dff06f", X"2006c583", X"00f50633", X"00178793", X"00b60023", X"fa9ff06f", X"100607b7",
        X"00300613", X"20c78423", X"fff00713", X"20e78023", X"00100693", X"20d78423", X"f9f00713", X"20e78023",
        X"2007c583", X"2007c703", X"20c78423", X"01f00793", X"0ff77713", X"02f59e63", X"02600793", X"02f71063",
        X"00d52423", X"000017b7", X"00f52623", X"00f52823", X"ff078793", X"00f52c23", X"00008067", X"02700793",
        X"00f71863", X"00d52423", X"000027b7", X"fddff06f", X"00000513", X"00008067", X"fe010113", X"000067b7",
        X"00812c23", X"00912a23", X"01212823", X"01312623", X"02c78793", X"00112e23", X"01412423", X"00f52023",
        X"8201c783", X"00050493", X"84c18413", X"04079463", X"01000513", X"00042223", X"4a5010ef", X"00a42023",
        X"00400513", X"499010ef", X"00400793", X"00a42423", X"00002537", X"00f42623", X"82818613", X"00100793",
        X"84c18593", X"54450513", X"00042823", X"82f18023", X"475010ef", X"01042a03", X"00c42783", X"06fa1263",
        X"01000913", X"000a0463", X"001a1913", X"01242623", X"200007b7", X"fff00513", X"00f97463", X"00291513",
        X"43d010ef", X"00050993", X"00090513", X"431010ef", X"00050913", X"00842683", X"00042503", X"00000793",
        X"0b47c463", X"00050463", X"419010ef", X"00842503", X"00050463", X"40d010ef", X"01342023", X"01242423",
        X"01042703", X"00042783", X"00271693", X"00d787b3", X"0097a023", X"00842783", X"00e787b3", X"00078023",
        X"01042783", X"01c12083", X"00a00713", X"00178793", X"00f42823", X"000067b7", X"0a878793", X"00f4a023",
        X"21000793", X"00f4a223", X"00100793", X"00f4a423", X"01812403", X"000017b7", X"00f4a623", X"00f4a823",
        X"ff078793", X"00e4aa23", X"00f4ac23", X"00048e23", X"01012903", X"01412483", X"00c12983", X"00812a03",
        X"02010113", X"00008067", X"00279713", X"00e50633", X"00062603", X"00e98733", X"00c72023", X"00f68733",
        X"00074603", X"00f90733", X"00178793", X"00c70023", X"f31ff06f", X"fe010113", X"00812c23", X"00912a23",
        X"01212823", X"01312623", X"00112e23", X"100607b7", X"00100713", X"20e78423", X"fd700713", X"20e78023",
        X"00050913", X"00058413", X"c10fd0ef", X"00050493", X"100609b7", X"2009c783", X"0ff7f793", X"00f90e23",
        X"01879793", X"4187d793", X"0207ce63", X"becfd0ef", X"409507b3", X"fef450e3", X"00000513", X"100607b7",
        X"00300713", X"20e78423", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"02010113",
        X"00008067", X"00100513", X"fd5ff06f", X"01852703", X"01452783", X"00e585b3", X"00f595b3", X"00100713",
        X"100607b7", X"20e78423", X"f8100713", X"20e78023", X"4105d713", X"0ff77713", X"20e78023", X"4085d713",
        X"0ff77713", X"20e78023", X"0ff5f593", X"20b78023", X"00300713", X"20e78423", X"1f400593", X"f19ff06f",
        X"01452783", X"fe010113", X"00812c23", X"00912a23", X"01312623", X"01412423", X"00112e23", X"01212823",
        X"01512223", X"00f595b3", X"00100693", X"100607b7", X"00452703", X"4105da13", X"20d78423", X"f8500693",
        X"20d78023", X"4085d993", X"0ffa7a13", X"21478023", X"0ff9f993", X"21378023", X"0ff5f413", X"20878023",
        X"00050493", X"40275713", X"00000793", X"100605b7", X"04e7c463", X"10060937", X"00300a93", X"21590423",
        X"1f400593", X"00048513", X"e8dff0ef", X"04051263", X"00000513", X"01c12083", X"01812403", X"01412483",
        X"01012903", X"00c12983", X"00812a03", X"00412a83", X"02010113", X"00008067", X"00279693", X"00d606b3",
        X"0006a683", X"00178793", X"20d5a023", X"fa5ff06f", X"00100793", X"20f90423", X"06100793", X"20f90023",
        X"21490023", X"21390023", X"20890023", X"21590423", X"1f400593", X"00048513", X"e1dff0ef", X"f8050ae3",
        X"01c4c503", X"00655513", X"00154513", X"00157513", X"f85ff06f", X"ff010113", X"00812423", X"00050413",
        X"00058513", X"00842583", X"00112623", X"565010ef", X"01442783", X"10060737", X"00100693", X"20d70423",
        X"00f517b3", X"07c00693", X"20d70023", X"4107d693", X"0ff6f693", X"20d70023", X"4087d693", X"0ff6f693",
        X"20d70023", X"0ff7f793", X"20f70023", X"00300793", X"20f70423", X"00040513", X"00812403", X"00c12083",
        X"000045b7", X"a9858593", X"01010113", X"d89ff06f", X"fe010113", X"00812c23", X"00912a23", X"01212823",
        X"01312623", X"00112e23", X"100604b7", X"00100993", X"3d2a8937", X"21348423", X"fcf90793", X"20f4a023",
        X"00300793", X"20f48423", X"06400593", X"00050413", X"d45ff0ef", X"08050063", X"21348423", X"00c42783",
        X"ffc90913", X"2124a023", X"4027d793", X"00179793", X"00000713", X"100606b7", X"fff00613", X"04f74063",
        X"100606b7", X"00c42703", X"04e7c063", X"100607b7", X"00300713", X"20e78423", X"00040513", X"01812403",
        X"01c12083", X"01412483", X"01012903", X"00c12983", X"06400593", X"02010113", X"cddff06f", X"20c68023",
        X"00170713", X"fb9ff06f", X"20068023", X"00178793", X"fb5ff06f", X"01c12083", X"01812403", X"01412483",
        X"01012903", X"00c12983", X"02010113", X"00008067", X"00c52503", X"00008067", X"00100513", X"00008067",
        X"00008067", X"100607b7", X"00100713", X"20e78423", X"00300713", X"20e78023", X"4105d713", X"0ff77713",
        X"20e78023", X"4085d713", X"0ff77713", X"20e78023", X"0ff5f593", X"20b78023", X"10060737", X"00000793",
        X"00c7ca63", X"100607b7", X"00300713", X"20e78423", X"00008067", X"20074503", X"00f685b3", X"00178793",
        X"00a58023", X"fddff06f", X"100606b7", X"00300593", X"20b68423", X"fff00713", X"20e68023", X"00100713",
        X"20e68423", X"f9f00713", X"20e68023", X"00050793", X"2006c503", X"2006c603", X"2006c703", X"20b68423",
        X"0ef00693", X"0ff67613", X"0ff77713", X"0ad51e63", X"04000693", X"00000513", X"0ad61a63", X"fec70713",
        X"0ff77713", X"00400693", X"0ae6e263", X"000066b7", X"00271713", X"18c68693", X"00d70733", X"00072703",
        X"00070067", X"01000713", X"00e7a223", X"10000713", X"00e7a423", X"00001737", X"00e7a623", X"00078513",
        X"00008067", X"01000713", X"00e7a223", X"20000713", X"00e7a423", X"00002737", X"fe1ff06f", X"01000713",
        X"00e7a223", X"40000713", X"00e7a423", X"00004737", X"fc9ff06f", X"01000713", X"00e7a223", X"00001737",
        X"80070713", X"00e7a423", X"00008737", X"fadff06f", X"01000713", X"00e7a223", X"00001737", X"00e7a423",
        X"00010737", X"f95ff06f", X"00000513", X"00008067", X"00c52783", X"00004737", X"04e78063", X"02f74063",
        X"00001737", X"04e78063", X"00002737", X"04e79863", X"00006537", X"1a850513", X"00008067", X"00008737",
        X"02e78863", X"00010737", X"02e79a63", X"00006537", X"1c050513", X"00008067", X"00006537", X"1b050513",
        X"00008067", X"00006537", X"1a050513", X"00008067", X"00006537", X"1b850513", X"00008067", X"00006537",
        X"1c850513", X"00008067", X"10000513", X"00008067", X"00052783", X"ff010113", X"00112623", X"0287a783",
        X"00812423", X"00050413", X"000780e7", X"00442583", X"201010ef", X"00c12083", X"00812403", X"01010113",
        X"00008067", X"00052783", X"01c7a783", X"00078067", X"100607b7", X"00100713", X"20e78423", X"04b00713",
        X"20e78023", X"2007a023", X"10060737", X"00000793", X"00800693", X"20074503", X"00f58633", X"00178793",
        X"00a60023", X"fed798e3", X"00300793", X"20f70423", X"00008067", X"00052783", X"ff010113", X"00112623",
        X"0287a783", X"000780e7", X"00c12083", X"00151513", X"01010113", X"00008067", X"01000513", X"00008067",
        X"00052783", X"fe010113", X"00112e23", X"04c7a783", X"00812c23", X"00912a23", X"01212823", X"00c12623",
        X"00d12423", X"00852903", X"00050413", X"00058493", X"000780e7", X"00442583", X"40a90533", X"00950533",
        X"131010ef", X"00042783", X"00851593", X"00040513", X"01812403", X"00812683", X"00c12603", X"01c12083",
        X"01412483", X"01012903", X"01c7a783", X"02010113", X"00078067", X"00052783", X"fe010113", X"00912a23",
        X"04c7a783", X"00852483", X"00112e23", X"00812c23", X"01212823", X"01312623", X"00050413", X"00060993",
        X"00058913", X"000780e7", X"00442583", X"40a484b3", X"012484b3", X"00048513", X"0b9010ef", X"00042783",
        X"00050913", X"00048593", X"0307a783", X"00040513", X"000780e7", X"00042783", X"00098613", X"00090593",
        X"0407a783", X"00040513", X"000780e7", X"00042783", X"00040513", X"0407a483", X"0287a783", X"000780e7",
        X"00a98633", X"00040513", X"01812403", X"01c12083", X"00c12983", X"00190593", X"00048793", X"01012903",
        X"01412483", X"02010113", X"00078067", X"00052783", X"ff010113", X"00812423", X"04c7a783", X"00912223",
        X"01212023", X"00112623", X"00050413", X"00058493", X"00852903", X"000780e7", X"00042783", X"40a905b3",
        X"00040513", X"00812403", X"00c12083", X"00012903", X"0307a783", X"009585b3", X"00412483", X"01010113",
        X"00078067", X"100607b7", X"00100713", X"20e78423", X"00859593", X"00300713", X"20e78023", X"4105d713",
        X"0ff77713", X"4085d593", X"20e78023", X"0ff5f593", X"20b78023", X"20078023", X"10060713", X"2007a683",
        X"00460613", X"fed62e23", X"fec71ae3", X"00300713", X"20e78423", X"00100513", X"00008067", X"ff010113",
        X"00812423", X"100607b7", X"00112623", X"00912223", X"01212023", X"20078423", X"00600713", X"20e78023",
        X"00100713", X"20e78423", X"00859593", X"00200713", X"20e78023", X"4105d713", X"0ff77713", X"4085d593",
        X"20e78023", X"0ff5f593", X"20b78023", X"20078023", X"10060437", X"10060793", X"00062703", X"00460613",
        X"20e42023", X"fec79ae3", X"00300493", X"20940423", X"00052783", X"00f00593", X"0707a783", X"000780e7",
        X"00400793", X"20040423", X"20f40023", X"20940423", X"00c12083", X"00812403", X"00412483", X"00012903",
        X"01010113", X"00008067", X"ff010113", X"00912223", X"00050493", X"00058513", X"0044a583", X"00112623",
        X"00812423", X"01212023", X"10060437", X"6c4010ef", X"00600713", X"20040423", X"20e40023", X"00100713",
        X"20e40423", X"00851793", X"02000713", X"20e40023", X"4107d713", X"0ff77713", X"4087d793", X"20e40023",
        X"0ff7f793", X"20f40023", X"20040023", X"00300913", X"21240423", X"0004a783", X"00048513", X"3e800593",
        X"0707a783", X"000780e7", X"00400793", X"20040423", X"20f40023", X"21240423", X"00c12083", X"00812403",
        X"00412483", X"00012903", X"01010113", X"00008067", X"00058793", X"00452583", X"ff010113", X"00078513",
        X"00112623", X"650010ef", X"00c12083", X"01010113", X"00008067", X"fd010113", X"02812423", X"00058413",
        X"000065b7", X"01400613", X"24c58593", X"00c10513", X"02112623", X"6ad010ef", X"01041713", X"01075713",
        X"00841793", X"00875713", X"00e7e7b3", X"00f11823", X"41045413", X"00300793", X"00f10a23", X"00810aa3",
        X"100607b7", X"60078223", X"60078223", X"10060737", X"00000793", X"01400693", X"00c10613", X"00f60633",
        X"00064603", X"00178793", X"60c70423", X"fed796e3", X"60070223", X"60070223", X"02c12083", X"02812403",
        X"03010113", X"00008067", X"fe010113", X"00112e23", X"00812c23", X"00912a23", X"01212823", X"01312623",
        X"01412423", X"10060437", X"20040423", X"00600a13", X"21440023", X"00100913", X"21240423", X"21240023",
        X"20040023", X"00300993", X"21340423", X"00052783", X"03200593", X"00050493", X"0707a783", X"000780e7",
        X"20040423", X"21440023", X"21240423", X"03100793", X"20f40023", X"20040023", X"21340423", X"0004a783",
        X"00048513", X"03200593", X"0707a783", X"000780e7", X"00400793", X"20040423", X"20f40023", X"01c12083",
        X"01812403", X"01412483", X"01012903", X"00c12983", X"00812a03", X"02010113", X"00008067", X"ff010113",
        X"00912223", X"100607b7", X"00112623", X"00812423", X"01212023", X"20078423", X"00600713", X"20e78023",
        X"00100713", X"20e78423", X"20e78023", X"00c52683", X"00008737", X"00050493", X"03800793", X"00e6c463",
        X"03400793", X"10060437", X"20f40023", X"00300913", X"21240423", X"0004a783", X"03200593", X"00048513",
        X"0707a783", X"000780e7", X"00600793", X"20040423", X"20f40023", X"00100793", X"20f40423", X"03100793",
        X"20f40023", X"20040023", X"21240423", X"0004a783", X"00048513", X"03200593", X"0707a783", X"000780e7",
        X"00400793", X"20040423", X"20f40023", X"00c12083", X"00812403", X"00412483", X"00012903", X"00100513",
        X"01010113", X"00008067", X"01000593", X"7cd0006f", X"ff010113", X"00812423", X"00912223", X"00112623",
        X"00058493", X"00060413", X"875fc0ef", X"040007b7", X"00f57533", X"04051c63", X"865fc0ef", X"020007b7",
        X"00f57533", X"04050a63", X"855fc0ef", X"300007b7", X"00f57533", X"04051863", X"000067b7", X"2c078593",
        X"0ff00713", X"0005c783", X"04e79463", X"00040513", X"01000613", X"44d010ef", X"00c12083", X"00812403",
        X"00412483", X"01010113", X"00008067", X"000067b7", X"31078593", X"fcdff06f", X"000067b7", X"26078593",
        X"fc1ff06f", X"000067b7", X"36078593", X"fb5ff06f", X"fa978ee3", X"01058593", X"fadff06f", X"fe010113",
        X"00812c23", X"00912a23", X"01212823", X"01312623", X"00112e23", X"00050493", X"00058413", X"00060993",
        X"00068913", X"fb8fc0ef", X"040007b7", X"00f57533", X"02051863", X"fa8fc0ef", X"020007b7", X"00f57533",
        X"02051663", X"000067b7", X"26078793", X"0ff00693", X"0007c703", X"02d71263", X"00000413", X"0480006f",
        X"000067b7", X"31078793", X"fe5ff06f", X"000067b7", X"2c078793", X"fd9ff06f", X"04871663", X"00c7a403",
        X"00895463", X"00090413", X"0004a703", X"0087a583", X"00098693", X"01c72703", X"00040613", X"00048513",
        X"000700e7", X"01c12083", X"00040513", X"01812403", X"01412483", X"01012903", X"00c12983", X"02010113",
        X"00008067", X"01078793", X"f89ff06f", X"ff010113", X"00812423", X"00912223", X"01212023", X"00112623",
        X"100607b7", X"00100713", X"20e78423", X"00500713", X"20e78023", X"00058493", X"f20fc0ef", X"00050413",
        X"10060937", X"20094783", X"0017f793", X"02079663", X"00100513", X"100607b7", X"00300713", X"20e78423",
        X"00c12083", X"00812403", X"00412483", X"00012903", X"01010113", X"00008067", X"ee0fc0ef", X"40850533",
        X"fca4d2e3", X"00000513", X"fcdff06f", X"100607b7", X"00100693", X"20d78423", X"00500693", X"20d78023",
        X"2007c683", X"00300613", X"20c78423", X"07c6f793", X"01000693", X"00d78863", X"00052783", X"0607a783",
        X"00078067", X"00008067", X"fe010113", X"000067b7", X"00812c23", X"00912a23", X"01212823", X"01312623",
        X"02c78793", X"00112e23", X"01412423", X"00f52023", X"8201c783", X"00050493", X"84c18413", X"04079463",
        X"01000513", X"00042223", X"555000ef", X"00a42023", X"00400513", X"549000ef", X"00400793", X"00a42423",
        X"00002537", X"00f42623", X"82818613", X"00100793", X"84c18593", X"54450513", X"00042823", X"82f18023",
        X"525000ef", X"01042a03", X"00c42783", X"06fa1263", X"01000913", X"000a0463", X"001a1913", X"01242623",
        X"200007b7", X"fff00513", X"00f97463", X"00291513", X"4ed000ef", X"00050993", X"00090513", X"4e1000ef",
        X"00050913", X"00842683", X"00042503", X"00000793", X"0947c863", X"00050463", X"4c9000ef", X"00842503",
        X"00050463", X"4bd000ef", X"01342023", X"01242423", X"01042703", X"00042783", X"00271693", X"00d787b3",
        X"0097a023", X"00842783", X"00e787b3", X"00078023", X"01042783", X"01c12083", X"01012903", X"00178793",
        X"00f42823", X"000067b7", X"1d878793", X"00f4a023", X"01000793", X"00f4a223", X"01812403", X"20000793",
        X"00f4a423", X"000027b7", X"00f4a623", X"00c12983", X"01412483", X"00812a03", X"02010113", X"00008067",
        X"00279713", X"00e50633", X"00062603", X"00e98733", X"00c72023", X"00f68733", X"00074603", X"00f90733",
        X"00178793", X"00c70023", X"f49ff06f", X"10060737", X"00050793", X"00300513", X"20a70423", X"fff00693",
        X"20d70023", X"00100593", X"20b70423", X"f9f00693", X"20d70023", X"20074803", X"20074603", X"20074683",
        X"20a70423", X"0ff67613", X"0ff6f693", X"04b81e63", X"04000713", X"00000513", X"04e61a63", X"01500713",
        X"02e69263", X"01000713", X"00e7a823", X"20000713", X"00e7aa23", X"00002737", X"00e7ac23", X"00078513",
        X"00008067", X"01600713", X"00000513", X"02e69063", X"01000713", X"00e7a823", X"40000713", X"00e7aa23",
        X"00004737", X"fd5ff06f", X"00000513", X"00008067", X"ff010113", X"00812423", X"00112623", X"10060437",
        X"20040423", X"00600793", X"20f40023", X"00100793", X"20f40423", X"20f40023", X"02000793", X"20f40023",
        X"20040023", X"00300793", X"20f40423", X"00052783", X"03200593", X"0707a783", X"000780e7", X"00400793",
        X"20040423", X"20f40023", X"00c12083", X"00812403", X"01010113", X"00008067", X"ff010113", X"00812423",
        X"00112623", X"10060437", X"20040423", X"00600793", X"20f40023", X"00100793", X"20f40423", X"20f40023",
        X"02800793", X"20f40023", X"20040023", X"00300793", X"20f40423", X"00052783", X"03200593", X"0707a783",
        X"000780e7", X"00400793", X"20040423", X"20f40023", X"00c12083", X"00812403", X"00100513", X"01010113",
        X"00008067", X"000067b7", X"3b878793", X"00f52023", X"ab0ff06f", X"ff010113", X"00812423", X"00112623",
        X"00050413", X"fe1ff0ef", X"00040513", X"00812403", X"00c12083", X"01c00593", X"01010113", X"25d0006f",
        X"100607b7", X"00100693", X"20d78423", X"00500693", X"20d78023", X"2007c683", X"00300613", X"20c78423",
        X"07c6f793", X"02800693", X"00d78863", X"00052783", X"0607a783", X"00078067", X"00008067", X"ff010113",
        X"00812423", X"00112623", X"00050413", X"c7dff0ef", X"000067b7", X"3b878793", X"00f42023", X"01000793",
        X"00f42823", X"20000793", X"00f42a23", X"000027b7", X"00c12083", X"00f42c23", X"00812403", X"01010113",
        X"00008067", X"ff010113", X"000067b7", X"00812423", X"00112623", X"64878793", X"00050413", X"00f52023",
        X"00006537", X"42c50513", X"cc1fd0ef", X"00040513", X"00812403", X"00c12083", X"01010113", X"d35fd06f",
        X"ff010113", X"00812423", X"00112623", X"00050413", X"fb5ff0ef", X"00040513", X"00812403", X"00c12083",
        X"01000593", X"01010113", X"1710006f", X"fe010113", X"00812c23", X"00112e23", X"00a12623", X"76c000ef",
        X"00157793", X"00c12583", X"00200413", X"00078663", X"00151793", X"0047f413", X"00d5c783", X"00079a63",
        X"00006537", X"45450513", X"bf5fd0ef", X"00146413", X"01c12083", X"00040513", X"01812403", X"02010113",
        X"00008067", X"00800793", X"100606b7", X"0ff00613", X"0006c703", X"0ff77513", X"00c71863", X"fff78793",
        X"0ff7f793", X"fe0796e3", X"00008067", X"ff010113", X"00812423", X"00112623", X"00050413", X"ca5fd0ef",
        X"000067b7", X"64878793", X"00c12083", X"00f42023", X"00042423", X"00041623", X"00812403", X"01010113",
        X"00008067", X"0ff00793", X"00f59863", X"00006537", X"47450513", X"bb5fd06f", X"ff010113", X"00812423",
        X"00112623", X"0405f793", X"00058413", X"00078863", X"00006537", X"48c50513", X"b91fd0ef", X"02047793",
        X"00078863", X"00006537", X"4a450513", X"b7dfd0ef", X"01047793", X"00078863", X"00006537", X"4bc50513",
        X"b69fd0ef", X"00847793", X"00078863", X"00006537", X"4dc50513", X"b55fd0ef", X"00447793", X"00078863",
        X"00006537", X"4e850513", X"b41fd0ef", X"00247793", X"00078863", X"00006537", X"4fc50513", X"b2dfd0ef",
        X"00147413", X"00040e63", X"00812403", X"00006537", X"00c12083", X"52450513", X"01010113", X"f59ff06f",
        X"00c12083", X"00812403", X"01010113", X"00008067", X"fe010113", X"00112e23", X"00812c23", X"01212823",
        X"01312623", X"00912a23", X"00052423", X"00051623", X"00050413", X"5e4000ef", X"0c800513", X"658000ef",
        X"06500913", X"00100993", X"00000613", X"00000593", X"00000513", X"5f8000ef", X"e8dff0ef", X"00050493",
        X"13350a63", X"fff90913", X"fe0910e3", X"0ff00793", X"00f50863", X"00048593", X"00040513", X"ec9ff0ef",
        X"00100493", X"01c12083", X"01812403", X"01012903", X"00c12983", X"00048513", X"01412483", X"02010113",
        X"00008067", X"00006537", X"53c50513", X"a5dfd0ef", X"00100793", X"00008937", X"00f42423", X"d0190913",
        X"00100993", X"00000613", X"00000593", X"03700513", X"57c000ef", X"e11ff0ef", X"000045b7", X"00000613",
        X"02900513", X"568000ef", X"dfdff0ef", X"00050593", X"00a9f863", X"00040513", X"e4dff0ef", X"f89ff06f",
        X"01351863", X"fff90913", X"fa091ee3", X"f75ff06f", X"00842703", X"00200793", X"04f71a63", X"00000613",
        X"00000593", X"03a00513", X"524000ef", X"db9ff0ef", X"00050593", X"00040513", X"e0dff0ef", X"100607b7",
        X"0007c703", X"fff00693", X"00d78023", X"00d78023", X"00d78023", X"04077793", X"00078a63", X"00006537",
        X"01340623", X"55050513", X"9a1fd0ef", X"00000513", X"524000ef", X"00006537", X"00040593", X"56050513",
        X"93dfd0ef", X"00100793", X"00f406a3", X"00000493", X"ef5ff06f", X"1aa00613", X"00000593", X"00800513",
        X"4ac000ef", X"d41ff0ef", X"00457513", X"ee051ce3", X"00006537", X"54450513", X"951fd0ef", X"100607b7",
        X"0007c703", X"fff00713", X"00e78023", X"0007c703", X"0007c703", X"0aa00793", X"eaf714e3", X"00200793",
        X"ed5ff06f", X"fe010113", X"00812c23", X"00912a23", X"01212823", X"01312623", X"01512223", X"00112e23",
        X"01412423", X"00050493", X"00058a93", X"00060413", X"00068993", X"00000913", X"00991a13", X"014a8a33",
        X"01394663", X"00000513", X"0400006f", X"00c4c783", X"00040593", X"00079463", X"00941593", X"01059613",
        X"01065613", X"0105d593", X"01100513", X"400000ef", X"c95ff0ef", X"00050593", X"02050a63", X"00048513",
        X"ce5ff0ef", X"00100513", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"00812a03",
        X"00412a83", X"02010113", X"00008067", X"000a0513", X"414000ef", X"00050593", X"fc0512e3", X"00140413",
        X"00190913", X"f75ff06f", X"fe010113", X"00812c23", X"00912a23", X"01212823", X"01312623", X"01512223",
        X"00112e23", X"01412423", X"00050913", X"00058a93", X"00060413", X"00068993", X"00000493", X"00949a13",
        X"014a8a33", X"0134c663", X"00000513", X"0580006f", X"00c94783", X"00040593", X"00079463", X"00941593",
        X"01059613", X"01065613", X"0105d593", X"01800513", X"33c000ef", X"bd1ff0ef", X"00050593", X"00090513",
        X"c25ff0ef", X"000a0513", X"40c000ef", X"02051e63", X"00006537", X"00040593", X"58450513", X"f80fd0ef",
        X"00100513", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"00812a03", X"00412a83",
        X"02010113", X"00008067", X"00140413", X"00148493", X"f6dff06f", X"fd010113", X"02912223", X"00000613",
        X"00058493", X"00a00513", X"00000593", X"02812423", X"03212023", X"02112623", X"01312e23", X"0c800413",
        X"2ac000ef", X"0fe00913", X"fff40413", X"b39ff0ef", X"0ff47413", X"01250c63", X"fe0418e3", X"00006537",
        X"61c50513", X"f44fd0ef", X"0600006f", X"fe0408e3", X"00000793", X"100605b7", X"01000713", X"0005c603",
        X"00f106b3", X"00178793", X"00c68023", X"fee798e3", X"00006537", X"61450513", X"ec4fd0ef", X"00000413",
        X"000069b7", X"01000913", X"008107b3", X"0007c583", X"5a498513", X"00140413", X"ea4fd0ef", X"ff2416e3",
        X"00a00513", X"f3cfd0ef", X"00000613", X"00000593", X"00900513", X"218000ef", X"0c800413", X"0fe00913",
        X"fff40413", X"aa1ff0ef", X"0ff47413", X"09250863", X"fe0418e3", X"100607b7", X"fff00713", X"00e78023",
        X"00e78023", X"0a040063", X"00006537", X"5ac50513", X"e4cfd0ef", X"00000413", X"000069b7", X"01000913",
        X"008107b3", X"0007c583", X"5a498513", X"00140413", X"e2cfd0ef", X"ff2416e3", X"00a00513", X"ec4fd0ef",
        X"00014683", X"00914783", X"00814703", X"0c06f693", X"08068463", X"00871713", X"00e787b3", X"01079413",
        X"01045413", X"00006537", X"00040593", X"5fc50513", X"decfd0ef", X"00a00913", X"0c00006f", X"f6040ce3",
        X"00000793", X"100605b7", X"01000713", X"0005c603", X"00f106b3", X"00178793", X"00c68023", X"fee798e3",
        X"f55ff06f", X"00006537", X"5b450513", X"dfcfd0ef", X"00000413", X"00100513", X"0084a023", X"02c12083",
        X"02812403", X"02412483", X"02012903", X"01c12983", X"03010113", X"00008067", X"00614403", X"00714683",
        X"00a14603", X"00347413", X"00269693", X"00675713", X"00e68733", X"00514583", X"00a41413", X"00e40433",
        X"00765613", X"00179793", X"01041413", X"00260613", X"0067f793", X"01045413", X"00f5f593", X"00f60633",
        X"00006537", X"00c58933", X"00040693", X"5c850513", X"ff790913", X"d28fd0ef", X"00140413", X"01241433",
        X"00000513", X"f75ff06f", X"00200713", X"04e58463", X"00b76863", X"02059c63", X"00000513", X"00008067",
        X"00300713", X"02e58e63", X"00006537", X"ff010113", X"63450513", X"00112623", X"ce4fd0ef", X"00c12083",
        X"00400513", X"01010113", X"00008067", X"00060593", X"d85ff06f", X"20000793", X"00f62023", X"fbdff06f",
        X"000207b7", X"ff5ff06f", X"100607b7", X"0087c503", X"00255513", X"00008067", X"100607b7", X"ffe00713",
        X"00e78223", X"00300713", X"00e78423", X"fff00693", X"06400793", X"10060737", X"00d70023", X"fff78793",
        X"fe079ce3", X"00070423", X"00008067", X"100607b7", X"fff00713", X"00e78023", X"00078623", X"04056513",
        X"00a78023", X"0085d713", X"00e78023", X"0ff5f593", X"00b78023", X"00865713", X"00e78023", X"0ff67613",
        X"00c78023", X"00c7c703", X"0ff77713", X"00e78023", X"00008067", X"0ff57513", X"100607b7", X"00a78223",
        X"00008067", X"0003b737", X"00050793", X"98070713", X"100605b7", X"0ff00613", X"0005c683", X"0ff6f513",
        X"04c68263", X"0fe00713", X"04e51263", X"0037f713", X"04071063", X"20078713", X"10060637", X"00062683",
        X"00478793", X"fed7ae23", X"fef71ae3", X"100607b7", X"fff00713", X"00e78023", X"00e78023", X"00000513",
        X"00c0006f", X"fff70713", X"fa0718e3", X"00008067", X"00000713", X"10060537", X"20000693", X"00054583",
        X"00e78633", X"00170713", X"00b60023", X"fed718e3", X"fbdff06f", X"100607b7", X"ffe00713", X"00e78023",
        X"00357793", X"04079863", X"20050793", X"10060737", X"00052683", X"00450513", X"00d72023", X"fea79ae3",
        X"100607b7", X"fff00713", X"00e78023", X"00e78023", X"00e78023", X"000927b7", X"7c078793", X"10060637",
        X"0ff00713", X"00064683", X"02e69863", X"00100513", X"00008067", X"00000793", X"100606b7", X"20000713",
        X"00f50633", X"00064603", X"00178793", X"00c68023", X"fee798e3", X"fadff06f", X"fff78793", X"fc0794e3",
        X"00000513", X"00008067", X"ff010113", X"00112623", X"538000ef", X"00051a63", X"00006537", X"66450513",
        X"b28fd0ef", X"0000006f", X"00c12083", X"01010113", X"00008067", X"fd5ff06f", X"5200006f", X"fcdff06f",
        X"5180006f", X"00008067", X"82a1ac23", X"00050067", X"fe010113", X"00c10613", X"00200593", X"00912a23",
        X"00112e23", X"00812c23", X"00050493", X"9c5fd0ef", X"00050e63", X"00000513", X"01c12083", X"01812403",
        X"01412483", X"02010113", X"00008067", X"00c12503", X"000017b7", X"e0078793", X"e0050713", X"fce7ece3",
        X"f9dff0ef", X"00050593", X"00050413", X"00100693", X"00000613", X"00048513", X"941fd0ef", X"00050593",
        X"00050a63", X"00006537", X"68c50513", X"a30fd0ef", X"fa5ff06f", X"1ff44783", X"1fe44703", X"00879793",
        X"00e7e7b3", X"0000b737", X"a5570713", X"f8e794e3", X"03744783", X"03644703", X"01000637", X"00879793",
        X"00e7e7b3", X"03844703", X"fff60613", X"005446b7", X"01071713", X"00f76733", X"03944783", X"14668693",
        X"00100513", X"01879793", X"00e7e7b3", X"00c7f7b3", X"f4d784e3", X"05344703", X"05244783", X"05544503",
        X"00871713", X"00f76733", X"05444783", X"01851513", X"01079793", X"00e7e7b3", X"00f56533", X"00c57533",
        X"40d50533", X"00153513", X"f11ff06f", X"ff010113", X"01800513", X"00112623", X"00812423", X"00912223",
        X"eb5ff0ef", X"8301a583", X"20000613", X"00050493", X"a84fd0ef", X"00000593", X"00048513", X"83418413",
        X"00942023", X"c94fd0ef", X"00050593", X"00050493", X"00006537", X"6cc50513", X"944fd0ef", X"fff00513",
        X"02905463", X"00042783", X"0147a403", X"00040513", X"e81ff0ef", X"02051463", X"00006537", X"6ec50513",
        X"968fd0ef", X"ffe00513", X"00c12083", X"00812403", X"00412483", X"01010113", X"00008067", X"8101c683",
        X"00069a63", X"00100693", X"80d18823", X"8081ac23", X"00c0006f", X"8181a703", X"fe070ae3", X"000065b7",
        X"00100613", X"70c58593", X"8bc18513", X"f68fc0ef", X"00050593", X"00050413", X"00006537", X"71050513",
        X"8bcfd0ef", X"00000513", X"fa0400e3", X"ffd00513", X"f99ff06f", X"ff010113", X"01000513", X"00112623",
        X"00812423", X"dd1ff0ef", X"00050413", X"ce0ff0ef", X"8281a823", X"00812403", X"00c12083", X"01010113",
        X"eedff06f", X"dc010113", X"22912a23", X"23212823", X"00100613", X"00050913", X"00058493", X"00050593",
        X"01010513", X"22812c23", X"22112e23", X"f70fc0ef", X"00050413", X"00050613", X"00006537", X"00090593",
        X"72850513", X"838fd0ef", X"04041463", X"00c10693", X"00400637", X"00048593", X"01010513", X"00012623",
        X"829fc0ef", X"00c12603", X"00006537", X"74450513", X"00060593", X"808fd0ef", X"01010513", X"a15fc0ef",
        X"00c12783", X"02078463", X"00048513", X"d3dff0ef", X"23c12083", X"00040513", X"23812403", X"23412483",
        X"23012903", X"24010113", X"00008067", X"00900413", X"fe1ff06f", X"fe010113", X"00112e23", X"00812c23",
        X"00912a23", X"01212823", X"891fd0ef", X"00052783", X"00010613", X"00200593", X"0207a783", X"00050413",
        X"000780e7", X"00042783", X"00812583", X"01c7a783", X"8ac18493", X"01000613", X"8ac18693", X"00040513",
        X"000780e7", X"0004c583", X"0014c783", X"00006537", X"01859593", X"01079793", X"00f5e5b3", X"0034c783",
        X"82c18913", X"00448613", X"00f5e5b3", X"0024c783", X"75c50513", X"00879793", X"00f5e5b3", X"00b92023",
        X"f3dfc0ef", X"00092603", X"fff00793", X"00000513", X"02f60663", X"00042783", X"00812583", X"000106b7",
        X"01c7a783", X"01058593", X"00040513", X"000780e7", X"00010537", X"c55ff0ef", X"00100513", X"01c12083",
        X"01812403", X"01412483", X"01012903", X"02010113", X"00008067", X"fe010113", X"004005b7", X"00010537",
        X"00112e23", X"decfb0ef", X"00050593", X"02055463", X"00a12623", X"00006537", X"78450513", X"ec1fc0ef",
        X"00c12583", X"01c12083", X"00058513", X"02010113", X"00008067", X"00006537", X"7a850513", X"ea1fc0ef",
        X"00010537", X"be5ff0ef", X"00100593", X"fd9ff06f", X"00050613", X"00000513", X"0015f693", X"00068463",
        X"00c50533", X"0015d593", X"00161613", X"fe0596e3", X"00008067", X"06054063", X"0605c663", X"00058613",
        X"00050593", X"fff00513", X"02060c63", X"00100693", X"00b67a63", X"00c05863", X"00161613", X"00169693",
        X"feb66ae3", X"00000513", X"00c5e663", X"40c585b3", X"00d56533", X"0016d693", X"00165613", X"fe0696e3",
        X"00008067", X"00008293", X"fb5ff0ef", X"00058513", X"00028067", X"40a00533", X"00b04863", X"40b005b3",
        X"f9dff06f", X"40b005b3", X"00008293", X"f91ff0ef", X"40a00533", X"00028067", X"00008293", X"0005ca63",
        X"00054c63", X"f79ff0ef", X"00058513", X"00028067", X"40b005b3", X"fe0558e3", X"40a00533", X"f61ff0ef",
        X"40b00533", X"00028067", X"000097b7", X"00050593", X"83c7a503", X"0140006f", X"000097b7", X"00050593",
        X"83c7a503", X"35d0006f", X"fd010113", X"01312e23", X"02112623", X"02812423", X"02912223", X"03212023",
        X"01412c23", X"01512a23", X"01612823", X"01712623", X"01812423", X"01912223", X"01a12023", X"00b58793",
        X"01600713", X"00050993", X"06f76663", X"01000793", X"1eb7e663", X"171000ef", X"01000493", X"01800793",
        X"00200613", X"00008937", X"00090913", X"00f907b3", X"0047a403", X"ff878713", X"20e40c63", X"00442783",
        X"00c42683", X"00842603", X"ffc7f793", X"00f407b3", X"0047a703", X"00d62623", X"00c6a423", X"00176713",
        X"00098513", X"00e7a223", X"121000ef", X"00840513", X"1980006f", X"ff87f493", X"1807c263", X"18b4e063",
        X"105000ef", X"1f700793", X"4697f663", X"0094d793", X"1a078863", X"00400713", X"3cf76c63", X"0064d793",
        X"03978613", X"03878513", X"00361693", X"00008937", X"00090913", X"00d906b3", X"0046a403", X"ff868693",
        X"02868663", X"00f00593", X"0100006f", X"32075c63", X"00c42403", X"00868c63", X"00442783", X"ffc7f793",
        X"40978733", X"fee5d4e3", X"00050613", X"01092403", X"00890893", X"17140a63", X"00442583", X"00f00713",
        X"ffc5f593", X"409587b3", X"40f74c63", X"01192a23", X"01192823", X"3e07d663", X"1ff00793", X"2eb7ea63",
        X"ff85f793", X"00878793", X"00492503", X"00f907b3", X"0007a683", X"0055d593", X"00100713", X"00b71733",
        X"00a76733", X"ff878593", X"00b42623", X"00d42423", X"00e92223", X"0087a023", X"0086a623", X"40265793",
        X"00100593", X"00f595b3", X"10b76a63", X"00e5f7b3", X"02079463", X"00159593", X"ffc67613", X"00e5f7b3",
        X"00460613", X"00079a63", X"00159593", X"00e5f7b3", X"00460613", X"fe078ae3", X"00f00813", X"00361313",
        X"00690333", X"00030513", X"00c52783", X"00060e13", X"2ef50263", X"0047a703", X"00078413", X"00c7a783",
        X"ffc77713", X"409706b3", X"2ed84263", X"fe06c2e3", X"00e40733", X"00472683", X"00842603", X"00098513",
        X"0016e693", X"00d72223", X"00f62623", X"00c7a423", X"798000ef", X"00840513", X"0100006f", X"00c00793",
        X"00f9a023", X"00000513", X"02c12083", X"02812403", X"02412483", X"02012903", X"01c12983", X"01812a03",
        X"01412a83", X"01012b03", X"00c12b83", X"00812c03", X"00412c83", X"00012d03", X"03010113", X"00008067",
        X"20000693", X"04000613", X"03f00513", X"e61ff06f", X"00c7a403", X"00260613", X"de8792e3", X"01092403",
        X"00890893", X"e9141ae3", X"00492703", X"40265793", X"00100593", X"00f595b3", X"eeb77ae3", X"00892403",
        X"00442b03", X"ffcb7b13", X"009b6863", X"409b07b3", X"00f00713", X"14f74463", X"00009c37", X"834c0c13",
        X"8441aa83", X"000c2703", X"fff00793", X"01640cb3", X"01548ab3", X"34f70863", X"000017b7", X"00f78793",
        X"00fa8ab3", X"fffff7b7", X"00fafab3", X"000a8593", X"00098513", X"6b8000ef", X"fff00793", X"00050b93",
        X"28f50a63", X"29956663", X"ae418d13", X"000d2a03", X"014a8a33", X"014d2023", X"000a0793", X"3aac8263",
        X"000c2683", X"fff00713", X"3ae68a63", X"419b8cb3", X"00fc87b3", X"00fd2023", X"007bfc13", X"300c0663",
        X"000017b7", X"418b8bb3", X"00878a13", X"008b8b93", X"418a0a33", X"015b8ab3", X"fff78793", X"415a0a33",
        X"00fa7a33", X"000a0593", X"00098513", X"640000ef", X"fff00793", X"3af50e63", X"41750533", X"01450ab3",
        X"000d2783", X"01792423", X"001aea93", X"00fa0a33", X"014d2023", X"015ba223", X"35240663", X"00f00693",
        X"3566f663", X"00442703", X"ff4b0793", X"ff87f793", X"00177713", X"00f76733", X"00e42223", X"00500613",
        X"00f40733", X"00c72223", X"00c72423", X"36f6ec63", X"004baa83", X"000b8413", X"83c18793", X"0007a703",
        X"01477463", X"0147a023", X"84018793", X"0007a703", X"1b477663", X"0147a023", X"1a40006f", X"0014e713",
        X"00e42223", X"009404b3", X"00992423", X"0017e793", X"00098513", X"00f4a223", X"590000ef", X"00840513",
        X"e09ff06f", X"00c42683", X"00842603", X"c41ff06f", X"0095d793", X"00400713", X"14f77263", X"01400713",
        X"22f76a63", X"05c78693", X"05b78713", X"00369693", X"00d906b3", X"0006a783", X"ff868693", X"1cf68863",
        X"0047a703", X"ffc77713", X"00e5f663", X"0087a783", X"fef698e3", X"00c7a683", X"00492703", X"00d42623",
        X"00f42423", X"0086a423", X"0087a623", X"cf1ff06f", X"01400713", X"12f77663", X"05400713", X"1ef76a63",
        X"00c4d793", X"06f78613", X"06e78513", X"00361693", X"c1dff06f", X"001e0e13", X"003e7793", X"00850513",
        X"10078e63", X"00c52783", X"d09ff06f", X"00842603", X"0014e593", X"00b42223", X"00f62623", X"00c7a423",
        X"009404b3", X"00992a23", X"00992823", X"0016e793", X"0114a623", X"0114a423", X"00f4a223", X"00e40733",
        X"00098513", X"00d72023", X"4a0000ef", X"00840513", X"d19ff06f", X"0034d613", X"00848793", X"b29ff06f",
        X"00b405b3", X"0045a783", X"00098513", X"0017e793", X"00f5a223", X"474000ef", X"00840513", X"cedff06f",
        X"0014e713", X"00e42223", X"009404b3", X"00992a23", X"00992823", X"0017e713", X"0114a623", X"0114a423",
        X"00e4a223", X"00b405b3", X"00098513", X"00f5a023", X"438000ef", X"00840513", X"cb1ff06f", X"0065d793",
        X"03978693", X"03878713", X"00369693", X"ec5ff06f", X"11240e63", X"00892403", X"00442a83", X"ffcafa93",
        X"409a87b3", X"009ae663", X"00f00713", X"e4f748e3", X"00098513", X"3f4000ef", X"00000513", X"c6dff06f",
        X"05c78613", X"05b78513", X"00361693", X"b01ff06f", X"00832783", X"fff60613", X"1c679063", X"00367793",
        X"ff830313", X"fe0796e3", X"00492703", X"fff5c793", X"00e7f7b3", X"00f92223", X"00159593", X"cab7e0e3",
        X"c8058ee3", X"00f5f733", X"00071a63", X"00159593", X"00f5f733", X"004e0e13", X"fe070ae3", X"000e0613",
        X"b9dff06f", X"010a8a93", X"cc5ff06f", X"00492503", X"40275593", X"00100713", X"00b71733", X"00a76733",
        X"00e92223", X"e39ff06f", X"015b8a33", X"41400a33", X"014a1a13", X"014a5a13", X"000a0593", X"00098513",
        X"34c000ef", X"fff00793", X"d0f518e3", X"00000a13", X"d11ff06f", X"05400713", X"08f76063", X"00c5d793",
        X"06f78693", X"06e78713", X"00369693", X"dc5ff06f", X"15400713", X"08f76063", X"00f4d793", X"07878613",
        X"07778513", X"00361693", X"a25ff06f", X"ae418d13", X"000d2783", X"00fa87b3", X"00fd2023", X"c65ff06f",
        X"014c9713", X"c4071ee3", X"00892403", X"015b0ab3", X"001aea93", X"01542223", X"d01ff06f", X"017c2023",
        X"c59ff06f", X"000b8413", X"cf1ff06f", X"00100793", X"00fba223", X"ebdff06f", X"15400713", X"06f76263",
        X"00f5d793", X"07878693", X"07778713", X"00369693", X"d41ff06f", X"55400713", X"06f76263", X"0124d793",
        X"07d78613", X"07c78513", X"00361693", X"9a1ff06f", X"ff8c0c13", X"018a8ab3", X"417a8ab3", X"00000a13",
        X"c41ff06f", X"00840593", X"00098513", X"3f4000ef", X"00892403", X"000d2a03", X"00442a83", X"c7dff06f",
        X"55400713", X"02f76463", X"0125d793", X"07d78693", X"07c78713", X"00369693", X"cd9ff06f", X"3f800693",
        X"07f00613", X"07e00513", X"945ff06f", X"3f800693", X"07e00713", X"cbdff06f", X"00492783", X"e5dff06f",
        X"00b547b3", X"0037f793", X"00c508b3", X"06079663", X"00300793", X"06c7f263", X"00357793", X"00050713",
        X"0c079a63", X"ffc8f613", X"40e606b3", X"02000793", X"02000293", X"06d7c263", X"00058693", X"00070793",
        X"02c77863", X"0006a803", X"00478793", X"00468693", X"ff07ae23", X"fec7e8e3", X"fff60793", X"40e787b3",
        X"ffc7f793", X"00478793", X"00f70733", X"00f585b3", X"01176863", X"00008067", X"00050713", X"ff157ce3",
        X"0005c783", X"00170713", X"00158593", X"fef70fa3", X"ff1768e3", X"00008067", X"0045a683", X"01c5a783",
        X"0005af83", X"0085af03", X"00c5ae83", X"0105ae03", X"0145a303", X"0185a803", X"00d72223", X"0205a683",
        X"01f72023", X"01e72423", X"01d72623", X"01c72823", X"00672a23", X"01072c23", X"00f72e23", X"02470713",
        X"40e607b3", X"fed72e23", X"02458593", X"faf2c6e3", X"f49ff06f", X"0005c683", X"00170713", X"00377793",
        X"fed70fa3", X"00158593", X"f0078ee3", X"0005c683", X"00170713", X"00377793", X"fed70fa3", X"00158593",
        X"fc079ae3", X"f01ff06f", X"00f00313", X"00050713", X"02c37e63", X"00f77793", X"0a079063", X"08059263",
        X"ff067693", X"00f67613", X"00e686b3", X"00b72023", X"00b72223", X"00b72423", X"00b72623", X"01070713",
        X"fed766e3", X"00061463", X"00008067", X"40c306b3", X"00269693", X"00000297", X"005686b3", X"00c68067",
        X"00b70723", X"00b706a3", X"00b70623", X"00b705a3", X"00b70523", X"00b704a3", X"00b70423", X"00b703a3",
        X"00b70323", X"00b702a3", X"00b70223", X"00b701a3", X"00b70123", X"00b700a3", X"00b70023", X"00008067",
        X"0ff5f593", X"00859693", X"00d5e5b3", X"01059693", X"00d5e5b3", X"f6dff06f", X"00279693", X"00000297",
        X"005686b3", X"00008293", X"fa0680e7", X"00028093", X"ff078793", X"40f70733", X"00f60633", X"f6c378e3",
        X"f3dff06f", X"00008067", X"00008067", X"ff010113", X"00812423", X"00912223", X"00050413", X"00058513",
        X"00112623", X"8401a423", X"e95fb0ef", X"fff00793", X"00f50c63", X"00c12083", X"00812403", X"00412483",
        X"01010113", X"00008067", X"8481a783", X"fe0784e3", X"00c12083", X"00f42023", X"00812403", X"00412483",
        X"01010113", X"00008067", X"fe010113", X"01312623", X"000089b7", X"00812c23", X"00912a23", X"01212823",
        X"01412423", X"00112e23", X"00058a13", X"00050913", X"00098993", X"f71ff0ef", X"0089a703", X"000017b7",
        X"fef78413", X"00472483", X"41440433", X"ffc4f493", X"00940433", X"00c45413", X"fff40413", X"00c41413",
        X"00f44e63", X"00000593", X"00090513", X"f41ff0ef", X"0089a783", X"009787b3", X"02f50863", X"00090513",
        X"f29ff0ef", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"00812a03", X"00000513",
        X"02010113", X"00008067", X"408005b3", X"00090513", X"efdff0ef", X"fff00793", X"04f50863", X"ae418793",
        X"0007a703", X"0089a683", X"408484b3", X"0014e493", X"40870733", X"00090513", X"0096a223", X"00e7a023",
        X"ec9ff0ef", X"01c12083", X"01812403", X"01412483", X"01012903", X"00c12983", X"00812a03", X"00100513",
        X"02010113", X"00008067", X"00000593", X"00090513", X"e9dff0ef", X"0089a703", X"00f00693", X"40e507b3",
        X"f4f6dee3", X"000096b7", X"8346a683", X"0017e793", X"00f72223", X"40d50533", X"aea1a223", X"f41ff06f",
        X"12058a63", X"ff010113", X"00812423", X"00912223", X"00058413", X"00050493", X"00112623", X"e49ff0ef",
        X"ffc42803", X"ff840713", X"000085b7", X"ffe87793", X"00f70633", X"00058593", X"00462683", X"0085a503",
        X"ffc6f693", X"1ac50a63", X"00d62223", X"00187813", X"00d60533", X"0a081063", X"ff842303", X"00452803",
        X"00008537", X"40670733", X"00872883", X"00850513", X"006787b3", X"00187813", X"14a88063", X"00c72303",
        X"0068a623", X"01132423", X"1e080263", X"0017e693", X"00d72223", X"00f62023", X"1ff00693", X"0af6e863",
        X"ff87f693", X"00868693", X"0045a503", X"00d586b3", X"0006a603", X"0057d813", X"00100793", X"010797b3",
        X"00a7e7b3", X"ff868513", X"00a72623", X"00c72423", X"00f5a223", X"00e6a023", X"00e62623", X"00812403",
        X"00c12083", X"00048513", X"00412483", X"01010113", X"d79ff06f", X"00452503", X"00157513", X"02051e63",
        X"00008537", X"00d787b3", X"00850513", X"00862683", X"0017e893", X"00f70833", X"16a68663", X"00c62603",
        X"00c6a623", X"00d62423", X"01172223", X"00f82023", X"f69ff06f", X"00008067", X"0017e693", X"fed42e23",
        X"00f62023", X"1ff00693", X"f4f6fce3", X"0097d693", X"00400613", X"0ed66a63", X"0067d693", X"03968813",
        X"03868613", X"00381813", X"01058833", X"00082683", X"ff880813", X"12d80663", X"0046a603", X"ffc67613",
        X"00c7f663", X"0086a683", X"fed818e3", X"00c6a803", X"01072623", X"00d72423", X"00812403", X"00c12083",
        X"00e82423", X"00048513", X"00412483", X"00e6a623", X"01010113", X"cb5ff06f", X"14081463", X"00c62583",
        X"00862603", X"00f686b3", X"00812403", X"00b62623", X"00c5a423", X"0016e793", X"00c12083", X"00f72223",
        X"00048513", X"00d70733", X"00412483", X"00d72023", X"01010113", X"c75ff06f", X"00187813", X"00d786b3",
        X"02081063", X"ff842503", X"40a70733", X"00c72783", X"00872603", X"00a686b3", X"00f62623", X"00c7a423",
        X"000097b7", X"0016e613", X"8387a783", X"00c72223", X"00e5a423", X"eaf6e4e3", X"8441a583", X"00048513",
        X"c89ff0ef", X"e99ff06f", X"01400613", X"02d67463", X"05400613", X"06d66463", X"00c7d693", X"06f68813",
        X"06e68613", X"00381813", X"f01ff06f", X"00d787b3", X"e9dff06f", X"05c68813", X"05b68613", X"00381813",
        X"ee9ff06f", X"00e5aa23", X"00e5a823", X"00a72623", X"00a72423", X"01172223", X"00f82023", X"e41ff06f",
        X"0045a503", X"40265613", X"00100793", X"00c797b3", X"00a7e7b3", X"00f5a223", X"ed9ff06f", X"15400613",
        X"00d66c63", X"00f7d693", X"07868813", X"07768613", X"00381813", X"e95ff06f", X"55400613", X"00d66c63",
        X"0127d693", X"07d68813", X"07c68613", X"00381813", X"e79ff06f", X"3f800813", X"07e00613", X"e6dff06f",
        X"0017e693", X"00d72223", X"00f62023", X"dd1ff06f", X"000001cc", X"00000200", X"00000234", X"3a783425",
        X"00000020", X"203a7025", X"00000000", X"78323025", X"00000020", X"00202020", X"00544146", X"33544146",
        X"00000032", X"2c2b2a22", X"3d3c3b3a", X"5d5b3f3e", X"00007f7c", X"41459a80", X"808f418e", X"49454545",
        X"8f8e4949", X"4f929290", X"55554f99", X"9b9a9959", X"9f9e9d9c", X"554f4941", X"a7a6a5a5", X"abaaa9a8",
        X"afaeadac", X"b3b2b1b0", X"b7b6b5b4", X"bbbab9b8", X"bfbebdbc", X"c3c2c1c0", X"c7c6c5c4", X"cbcac9c8",
        X"cfcecdcc", X"d3d2d1d0", X"d7d6d5d4", X"dbdad9d8", X"dfdedddc", X"e3e2e1e0", X"e7e6e5e4", X"ebeae9e8",
        X"efeeedec", X"f3f2f1f0", X"f7f6f5f4", X"fbfaf9f8", X"fffefdfc", X"6c756e28", X"0000296c", X"00001c1c",
        X"00001bb4", X"00001a40", X"000019b4", X"000019b4", X"000019b4", X"000019b4", X"00001a40", X"000019b4",
        X"000019b4", X"000019b4", X"000019b4", X"000019b4", X"000019b4", X"00001bd0", X"000019b4", X"000019b4",
        X"00001b68", X"000019b4", X"00001a40", X"000019b4", X"000019b4", X"00001bf4", X"33323130", X"37363534",
        X"42413938", X"46454443", X"00000000", X"00000000", X"00000000", X"00001df0", X"00001e18", X"00001df4",
        X"00001e00", X"00001e08", X"00001e08", X"00001e10", X"20524245", X"72617453", X"25203a74", X"69532064",
        X"203a657a", X"54206425", X"3a657079", X"0a642520", X"00000000", X"75746552", X"6e696e72", X"20312067",
        X"74726170", X"6f697469", X"0000006e", X"6e696f47", X"6f742067", X"61657220", X"61702064", X"74697472",
        X"206e6f69", X"6c626174", X"70202e65", X"69747261", X"6e6f6974", X"73696c5f", X"73692074", X"0a702520",
        X"00000000", X"2052424d", X"72617453", X"25203a74", X"69532064", X"203a657a", X"54206425", X"3a657079",
        X"0a642520", X"00000000", X"75736552", X"6f20746c", X"42452066", X"65722052", X"203a6461", X"0a2e6425",
        X"00000000", X"74726150", X"6f697469", X"7263206e", X"65746165", X"25202164", X"00000a70", X"65736142",
        X"00000000", X"00000000", X"00000000", X"00002484", X"00002588", X"00002488", X"00002490", X"0000249c",
        X"000024a0", X"000024a8", X"000024ac", X"000024b0", X"000024b4", X"000024bc", X"000024c4", X"000024cc",
        X"000024d4", X"000024dc", X"000024e4", X"000024f0", X"000024f8", X"00002500", X"00002508", X"00002510",
        X"00002524", X"00002528", X"0000252c", X"00002530", X"00002538", X"0000253c", X"00002540", X"00206225",
        X"00000000", X"00000000", X"00002778", X"00002b20", X"00002cfc", X"00002490", X"00002930", X"0000284c",
        X"000028b8", X"000027c0", X"0000277c", X"00002768", X"00002824", X"0000282c", X"00003114", X"00002ab4",
        X"000029d8", X"00002a54", X"00003000", X"00002770", X"00002994", X"000029a0", X"000029a8", X"000029c4",
        X"00002fac", X"00002b28", X"00003190", X"00002ad8", X"00002afc", X"00002c20", X"613299aa", X"81320000",
        X"a1320000", X"a1304f00", X"00200e00", X"00000100", X"00000000", X"00000000", X"00053ca0", X"00000101",
        X"00053ca0", X"000a2800", X"0000e2e0", X"00000102", X"00061f80", X"000be000", X"000c6000", X"000000fd",
        X"00127f80", X"0023e000", X"000df000", X"000000fe", X"0020df00", X"003fc000", X"00002100", X"000000ff",
        X"0020dcf0", X"003fbc00", X"00000210", X"00003364", X"00003384", X"0000339c", X"000033b4", X"000033d0",
        X"51353257", X"00003038", X"51353257", X"00003631", X"51353257", X"00003233", X"51353257", X"00003436",
        X"51353257", X"00383231", X"626e6957", X"00646e6f", X"00000000", X"00000000", X"00003280", X"00003a88",
        X"000032e8", X"000033f0", X"000034b0", X"00003b3c", X"000034a4", X"00003284", X"00003a90", X"00003270",
        X"00003468", X"00003470", X"000037a8", X"00003850", X"000036a4", X"000024e4", X"000036fc", X"00003278",
        X"000034f4", X"00003518", X"00003520", X"00003594", X"0000364c", X"00003874", X"000039bc", X"00003908",
        X"00003c8c", X"00002540", X"00003c0c", X"613299aa", X"81320000", X"a1320000", X"a1304f00", X"00200e00",
        X"00000100", X"00000000", X"00000000", X"00053ca0", X"00000101", X"00054000", X"00054000", X"0000e000",
        X"00000102", X"00062000", X"00062000", X"000c6000", X"000000fd", X"00128000", X"00128000", X"000c8000",
        X"000000fe", X"001f0000", X"001f0000", X"00010000", X"000000ff", X"001fe000", X"001fe000", X"00001000",
        X"00000000", X"00000000", X"00000000", X"000c0000", X"00000002", X"000c0000", X"000c0000", X"00140000",
        X"000000fd", X"00200000", X"00200000", X"001f0000", X"000000fe", X"003f0000", X"003f0000", X"00010000",
        X"000000ff", X"003fe000", X"003fe000", X"00001000", X"00000000", X"00000000", X"00000000", X"00290000",
        X"00000002", X"00290000", X"00290000", X"00170000", X"000000fd", X"00400000", X"00400000", X"003e8000",
        X"000000fe", X"007e8000", X"007e8000", X"00018000", X"000000ff", X"007fe000", X"007fe000", X"00001000",
        X"00000000", X"00000000", X"00000000", X"000c0000", X"00000002", X"000a0000", X"000a0000", X"00160000",
        X"000000fd", X"00200000", X"00200000", X"005f0000", X"000000fe", X"007f0000", X"007f0000", X"00010000",
        X"000000ff", X"007fe000", X"007fe000", X"00001000", X"00000000", X"00000000", X"00003fc4", X"00003fd4",
        X"00003e4c", X"000033f0", X"000034b0", X"00003b3c", X"000034a4", X"00003284", X"00003a90", X"00003270",
        X"00003468", X"00003470", X"000037a8", X"00003850", X"000036a4", X"000024e4", X"000036fc", X"00003278",
        X"000034f4", X"00003518", X"00003520", X"00003594", X"0000364c", X"00003874", X"00003f58", X"00003ef0",
        X"00004000", X"00002540", X"00003c0c", X"44202a2a", X"52545345", X"49544355", X"5320474e", X"52414344",
        X"4c422044", X"444b434f", X"43495645", X"2a2a2045", X"00000000", X"61436453", X"6e206472", X"6920746f",
        X"6974696e", X"7a696c61", X"2e2e6465", X"0a702520", X"00000000", X"78656e55", X"74636570", X"49206465",
        X"20454c44", X"65747962", X"0000002e", X"75677241", X"746e656d", X"74756f20", X"20666f20", X"6e756f62",
        X"002e7364", X"72646441", X"20737365", X"2074756f", X"6220666f", X"646e756f", X"00002e73", X"6f727245",
        X"75642072", X"676e6972", X"61726520", X"73206573", X"65757165", X"2e65636e", X"00000000", X"20435243",
        X"6c696166", X"002e6465", X"656c6c49", X"206c6167", X"6d6d6f63", X"2e646e61", X"00000000", X"73617245",
        X"65722065", X"20746573", X"65657328", X"6e615320", X"6b736944", X"636f6420", X"35702073", X"2933312d",
        X"0000002e", X"64726143", X"20736920", X"74696e69", X"696c6169", X"676e6973", X"0000002e", X"56204453",
        X"00782e31", X"56204453", X"30302e32", X"00000000", X"68676948", X"70616320", X"74696361", X"00002179",
        X"74746553", X"20676e69", X"74696e69", X"696c6169", X"2064657a", X"74206f74", X"2e657572", X"7025202e",
        X"0000000a", X"656d6954", X"2074756f", X"6f727265", X"72772072", X"6e697469", X"6c622067", X"206b636f",
        X"000a6425", X"32302520", X"00000078", X"3a445343", X"00000000", X"6c696146", X"74206465", X"6572206f",
        X"43206461", X"002e4453", X"64616572", X"5f6c625f", X"65776f70", X"203d2072", X"202e6425", X"657a6973",
        X"776f705f", X"3d207265", X"2e642520", X"735f6320", X"20657a69", X"6425203d", X"00000a2e", X"20445343",
        X"3a302e32", X"735f6320", X"20657a69", X"6425203d", X"00000a2e", X"3a444943", X"00000020", X"6c696146",
        X"74206465", X"6572206f", X"43206461", X"20647261", X"002e4449", X"54434f49", X"6425204c", X"00000a2e",
        X"00000000", X"00000000", X"00004084", X"000040c0", X"00004270", X"000040ec", X"00004444", X"00004508",
        X"00004808", X"50202a2a", X"43494e41", X"3a2a2a20", X"72724520", X"6120726f", X"636f6c6c", X"6e697461",
        X"656d2067", X"79726f6d", X"00002e2e", X"656c6946", X"74737953", X"41466d65", X"743a3a54", X"20747365",
        X"6c696166", X"202c6465", X"61636562", X"20657375", X"64616572", X"20676e69", X"74636573", X"6620726f",
        X"656c6961", X"25203a64", X"00000a64", X"6b736944", X"696e6920", X"6c616974", X"64657a69", X"6552202e",
        X"6e727574", X"203a6465", X"000a6425", X"20646944", X"20746f6e", X"646e6966", X"54414620", X"6c696620",
        X"79732065", X"6d657473", X"0000002e", X"00003a30", X"6e756f4d", X"20534674", X"75746572", X"64656e72",
        X"6425203a", X"0000000a", X"656c6946", X"20732520", X"6e65706f", X"73657220", X"20746c75", X"6425203d",
        X"00000a2e", X"65747942", X"65722073", X"203a6461", X"28206425", X"36257830", X"000a2978", X"6c707041",
        X"74616369", X"206e6f69", X"676e656c", X"3d206874", X"38302520", X"76202c78", X"69737265", X"25206e6f",
        X"00000a73", X"646f6d58", X"72206d65", X"69656365", X"65206576", X"726f7272", X"7473203a", X"73757461",
        X"6425203a", X"0000000a", X"646f6d58", X"73206d65", X"65636375", X"75667373", X"20796c6c", X"65636572",
        X"64657669", X"20642520", X"65747962", X"00000a73", X"322e3356", X"00000000", X"202a2a2a", X"31343531",
        X"746c5520", X"74616d69", X"49492d65", X"42202d20", X"6c746f6f", X"6564616f", X"73252072", X"46202d20",
        X"20414750", X"73726556", X"3a6e6f69", X"78322520", X"2a2a2a20", X"00000a0a", X"61647075", X"752e6574",
        X"00007232", X"69746c75", X"6574616d", X"6e69622e", X"00000000", X"656c6946", X"73797320", X"206d6574",
        X"6f727265", X"25203a72", X"00000a64", X"756f590a", X"20657227", X"64616564", X"00000021", X"00000000",
        X"00000000", X"00008000", X"00008000", X"00008008", X"00008008", X"00008010", X"00008010", X"00008018",
        X"00008018", X"00008020", X"00008020", X"00008028", X"00008028", X"00008030", X"00008030", X"00008038",
        X"00008038", X"00008040", X"00008040", X"00008048", X"00008048", X"00008050", X"00008050", X"00008058",
        X"00008058", X"00008060", X"00008060", X"00008068", X"00008068", X"00008070", X"00008070", X"00008078",
        X"00008078", X"00008080", X"00008080", X"00008088", X"00008088", X"00008090", X"00008090", X"00008098",
        X"00008098", X"000080a0", X"000080a0", X"000080a8", X"000080a8", X"000080b0", X"000080b0", X"000080b8",
        X"000080b8", X"000080c0", X"000080c0", X"000080c8", X"000080c8", X"000080d0", X"000080d0", X"000080d8",
        X"000080d8", X"000080e0", X"000080e0", X"000080e8", X"000080e8", X"000080f0", X"000080f0", X"000080f8",
        X"000080f8", X"00008100", X"00008100", X"00008108", X"00008108", X"00008110", X"00008110", X"00008118",
        X"00008118", X"00008120", X"00008120", X"00008128", X"00008128", X"00008130", X"00008130", X"00008138",
        X"00008138", X"00008140", X"00008140", X"00008148", X"00008148", X"00008150", X"00008150", X"00008158",
        X"00008158", X"00008160", X"00008160", X"00008168", X"00008168", X"00008170", X"00008170", X"00008178",
        X"00008178", X"00008180", X"00008180", X"00008188", X"00008188", X"00008190", X"00008190", X"00008198",
        X"00008198", X"000081a0", X"000081a0", X"000081a8", X"000081a8", X"000081b0", X"000081b0", X"000081b8",
        X"000081b8", X"000081c0", X"000081c0", X"000081c8", X"000081c8", X"000081d0", X"000081d0", X"000081d8",
        X"000081d8", X"000081e0", X"000081e0", X"000081e8", X"000081e8", X"000081f0", X"000081f0", X"000081f8",
        X"000081f8", X"00008200", X"00008200", X"00008208", X"00008208", X"00008210", X"00008210", X"00008218",
        X"00008218", X"00008220", X"00008220", X"00008228", X"00008228", X"00008230", X"00008230", X"00008238",
        X"00008238", X"00008240", X"00008240", X"00008248", X"00008248", X"00008250", X"00008250", X"00008258",
        X"00008258", X"00008260", X"00008260", X"00008268", X"00008268", X"00008270", X"00008270", X"00008278",
        X"00008278", X"00008280", X"00008280", X"00008288", X"00008288", X"00008290", X"00008290", X"00008298",
        X"00008298", X"000082a0", X"000082a0", X"000082a8", X"000082a8", X"000082b0", X"000082b0", X"000082b8",
        X"000082b8", X"000082c0", X"000082c0", X"000082c8", X"000082c8", X"000082d0", X"000082d0", X"000082d8",
        X"000082d8", X"000082e0", X"000082e0", X"000082e8", X"000082e8", X"000082f0", X"000082f0", X"000082f8",
        X"000082f8", X"00008300", X"00008300", X"00008308", X"00008308", X"00008310", X"00008310", X"00008318",
        X"00008318", X"00008320", X"00008320", X"00008328", X"00008328", X"00008330", X"00008330", X"00008338",
        X"00008338", X"00008340", X"00008340", X"00008348", X"00008348", X"00008350", X"00008350", X"00008358",
        X"00008358", X"00008360", X"00008360", X"00008368", X"00008368", X"00008370", X"00008370", X"00008378",
        X"00008378", X"00008380", X"00008380", X"00008388", X"00008388", X"00008390", X"00008390", X"00008398",
        X"00008398", X"000083a0", X"000083a0", X"000083a8", X"000083a8", X"000083b0", X"000083b0", X"000083b8",
        X"000083b8", X"000083c0", X"000083c0", X"000083c8", X"000083c8", X"000083d0", X"000083d0", X"000083d8",
        X"000083d8", X"000083e0", X"000083e0", X"000083e8", X"000083e8", X"000083f0", X"000083f0", X"000083f8",
        X"000083f8", X"00000000", X"000086f4", X"0000875c", X"000087c4", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000001", X"00000000", X"abcd330e", X"e66d1234", X"0005deec",
        X"0000000b", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00008b4c", X"ffffffff", X"00020000", X"00008408", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000"

    );
end package;
