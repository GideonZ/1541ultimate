
library ieee;
use ieee.std_logic_1164.all;

package bootrom_pkg is
    type t_boot_data    is array(natural range <>) of std_logic_vector(31 downto 0);

    constant c_bootrom : t_boot_data(0 to 2047) := (
        X"30047073", X"00002117", X"ff810113", X"00002197", X"3f418193", X"00000517", X"0cc50513", X"30551073",
        X"34151073", X"30001073", X"30401073", X"34401073", X"32001073", X"30601073", X"b0001073", X"b8001073",
        X"b0201073", X"b8201073", X"00000093", X"00000213", X"00000293", X"00000313", X"00000393", X"00001597",
        X"d8058593", X"00002617", X"b9c60613", X"00002697", X"b9468693", X"00d65c63", X"0005a703", X"00e62023",
        X"00458593", X"00460613", X"fedff06f", X"00002717", X"b7470713", X"80818793", X"00f75863", X"00072023",
        X"00470713", X"ff5ff06f", X"00000513", X"00000593", X"088000ef", X"34051073", X"10500073", X"0000006f",
        X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013", X"00000013",
        X"ff810113", X"00812023", X"00912223", X"34202473", X"02044663", X"34102473", X"00041483", X"0034f493",
        X"00240413", X"34141073", X"00300413", X"00941863", X"34102473", X"00240413", X"34141073", X"10000437",
        X"04900493", X"00940fa3", X"00012403", X"00412483", X"00810113", X"30200073", X"80001537", X"fe010113",
        X"d0c50513", X"00812c23", X"00112e23", X"00912a23", X"01212823", X"01312623", X"01412423", X"01512223",
        X"1cd000ef", X"bfc1a783", X"0007a783", X"02079063", X"000095b7", X"10058593", X"00000513", X"2ad000ef",
        X"bfc1a783", X"00100713", X"00e7a023", X"10060437", X"00300a13", X"21440423", X"fff00993", X"21340023",
        X"00100a93", X"21540423", X"21340023", X"21440423", X"1d5000ef", X"00050493", X"10100937", X"404000ef",
        X"00c94503", X"174000ef", X"0404d863", X"1b8000ef", X"1571c4b7", X"00010437", X"abe48493", X"800019b7",
        X"80001a37", X"ffc42783", X"14979263", X"d7898513", X"41c000ef", X"fe042e23", X"ff842903", X"00090513",
        X"3c0000ef", X"d4ca0513", X"404000ef", X"00090513", X"124000ef", X"fd1ff06f", X"70090423", X"488000ef",
        X"00010937", X"160000ef", X"ffc92703", X"1571c7b7", X"abe78793", X"02f71663", X"80001537", X"d2450513",
        X"3cc000ef", X"fe092e23", X"ff892503", X"0e8000ef", X"80001537", X"d5050513", X"3b4000ef", X"f75ff06f",
        X"400007b7", X"00f4f4b3", X"fe0494e3", X"21540423", X"21440023", X"02200793", X"20f40023", X"20040023",
        X"20040023", X"20042903", X"20042483", X"20042403", X"00090513", X"32c000ef", X"00048513", X"324000ef",
        X"00040513", X"31c000ef", X"80001537", X"d2c50513", X"35c000ef", X"f9348ee3", X"001807b7", X"00090513",
        X"fff48493", X"ffe78793", X"10060737", X"0297fe63", X"100607b7", X"80001537", X"20078423", X"d3c50513",
        X"32c000ef", X"100007b7", X"00a7c783", X"0077d793", X"02079663", X"00040513", X"03c000ef", X"00000013",
        X"00000013", X"ff9ff06f", X"20072683", X"ffc48493", X"00450513", X"fed52e23", X"fb5ff06f", X"80001537",
        X"d4850513", X"2e8000ef", X"fd5ff06f", X"00000013", X"eb5ff06f", X"00050067", X"ff010113", X"00812423",
        X"80001437", X"d8040413", X"00455793", X"00f407b3", X"00912223", X"00050493", X"0007c503", X"00f4f493",
        X"00112623", X"00940433", X"04d000ef", X"00044503", X"00812403", X"00c12083", X"00412483", X"01010113",
        X"0350006f", X"030307b7", X"fe010113", X"05778793", X"00f12023", X"0822d7b7", X"00278793", X"00f12223",
        X"010107b7", X"05778793", X"00f12423", X"8982f7b7", X"75578793", X"00912a23", X"101004b7", X"00812c23",
        X"00f12623", X"00112e23", X"7074c503", X"70048413", X"f69ff0ef", X"00a00513", X"7dc000ef", X"00c4c783",
        X"0037d793", X"feb78793", X"00f03733", X"00e40323", X"fc800713", X"70e48023", X"00144703", X"01871713",
        X"41875713", X"16074663", X"01400713", X"00e40023", X"10100737", X"70070713", X"00174683", X"01869693",
        X"4186d693", X"1406ca63", X"00800693", X"00d70023", X"101006b7", X"70068693", X"0016c703", X"01871713",
        X"41875713", X"12074e63", X"00000713", X"101005b7", X"00800513", X"00e106b3", X"0006c683", X"70058613",
        X"70d58023", X"00164683", X"01869693", X"4186d693", X"1006cc63", X"00170713", X"fca71ee3", X"00100713",
        X"00e601a3", X"10100737", X"70070713", X"00174683", X"01869693", X"4186d693", X"0e06cc63", X"0017b793",
        X"00f70323", X"fc800793", X"00f70023", X"101007b7", X"70078793", X"0017c703", X"01871713", X"41875713",
        X"0c074c63", X"01400713", X"00e78023", X"101007b7", X"70078793", X"0017c703", X"01871713", X"41875713",
        X"0c074063", X"00800713", X"00e78023", X"10100737", X"70070713", X"00174783", X"01879793", X"4187d793",
        X"0a07c463", X"00000793", X"10100637", X"00800593", X"00810713", X"00f70733", X"00074703", X"70060693",
        X"70e60023", X"0016c703", X"01871713", X"41875713", X"08074063", X"00178793", X"fcb79ce3", X"00100793",
        X"10100737", X"00f681a3", X"70070713", X"00174783", X"01879793", X"4187d793", X"0607c063", X"01c12083",
        X"01812403", X"01412483", X"02010113", X"00008067", X"00000013", X"e85ff06f", X"00000013", X"e9dff06f",
        X"00000013", X"eb5ff06f", X"00000013", X"ed9ff06f", X"00000013", X"ef9ff06f", X"00000013", X"f19ff06f",
        X"00000013", X"f31ff06f", X"00000013", X"f49ff06f", X"00000013", X"f71ff06f", X"00000013", X"f91ff06f",
        X"ff010113", X"00812423", X"00050413", X"01855513", X"00112623", X"d65ff0ef", X"01045513", X"0ff57513",
        X"d59ff0ef", X"00845513", X"0ff57513", X"d4dff0ef", X"0ff47513", X"d45ff0ef", X"00812403", X"00c12083",
        X"02000513", X"01010113", X"5ac0006f", X"ff010113", X"00812423", X"00112623", X"00050413", X"00044503",
        X"00051a63", X"00c12083", X"00812403", X"01010113", X"00008067", X"00140413", X"57c000ef", X"fe1ff06f",
        X"101007b7", X"10078713", X"10a79023", X"00b70123", X"00a00793", X"00274683", X"fff78793", X"fe079ce3",
        X"00008067", X"ff010113", X"00812423", X"00050413", X"00855513", X"00112623", X"00912223", X"00058493",
        X"cb9ff0ef", X"0ff47513", X"cb1ff0ef", X"00812403", X"00c12083", X"00048513", X"00412483", X"01010113",
        X"48c0006f", X"f4010113", X"0a912a23", X"101004b7", X"0a812c23", X"0a112e23", X"0b212823", X"0b312623",
        X"0b412423", X"0b512223", X"0b612023", X"09712e23", X"09812c23", X"09912a23", X"10048493", X"00900793",
        X"00f48623", X"7d000413", X"00c4c783", X"fff40413", X"fe041ce3", X"00200593", X"40000513", X"f45ff0ef",
        X"00000593", X"0000c537", X"f39ff0ef", X"00000593", X"00008537", X"f2dff0ef", X"00004537", X"00000593",
        X"05a50513", X"f1dff0ef", X"00000593", X"74200513", X"f11ff0ef", X"00200593", X"40000513", X"f05ff0ef",
        X"00100593", X"40000513", X"ef9ff0ef", X"00100593", X"40000513", X"eedff0ef", X"00100593", X"40000513",
        X"ee1ff0ef", X"00100593", X"40000513", X"ed5ff0ef", X"101007b7", X"00c7c783", X"01500713", X"0037d793",
        X"00e79663", X"00100793", X"00f484a3", X"123457b7", X"67878793", X"10f02023", X"876547b7", X"32178793",
        X"10f02223", X"00100713", X"101007b7", X"10e781a3", X"00a00513", X"400000ef", X"00000a93", X"fff00c93",
        X"05500b93", X"101006b7", X"01010793", X"10068713", X"00300613", X"10002583", X"00478793", X"00b12623",
        X"1046a583", X"feb7ae23", X"00c70323", X"01970223", X"019702a3", X"09010593", X"fcf59ee3", X"00000493",
        X"01f00b13", X"02000c13", X"01010793", X"00f48533", X"fff00a13", X"fff00913", X"00000613", X"00000793",
        X"02fb5c63", X"09991663", X"00148493", X"00400793", X"fcf49ce3", X"101007b7", X"00100713", X"10e783a3",
        X"001a8a93", X"f89a90e3", X"80001537", X"d9450513", X"2dc000ef", X"1400006f", X"00279713", X"00e50733",
        X"00074703", X"00178693", X"01770663", X"00068793", X"fb1ff06f", X"00078713", X"00070593", X"00170713",
        X"01870a63", X"00271693", X"00d506b3", X"0006c683", X"ff7684e3", X"40f586b3", X"00d65863", X"00058a13",
        X"00078913", X"00068613", X"00070793", X"f75ff06f", X"04600513", X"300000ef", X"0ff97513", X"a7dff0ef",
        X"04c00513", X"2f0000ef", X"0ffa7513", X"a6dff0ef", X"02091663", X"00900793", X"ff7a0993", X"0347c863",
        X"412a07b3", X"00a00713", X"fff00993", X"02f75063", X"014909b3", X"4019d993", X"0140006f", X"ff6a12e3",
        X"01600793", X"00990993", X"fd27cce3", X"04300513", X"2a4000ef", X"0ff9f913", X"00090513", X"a1dff0ef",
        X"00a00513", X"290000ef", X"f13050e3", X"101007b7", X"0ff4f493", X"10078793", X"00000713", X"00300613",
        X"fff00693", X"00978423", X"00c78323", X"00d78223", X"00d782a3", X"00170713", X"ff3748e3", X"04200513",
        X"254000ef", X"0ffaf513", X"9d1ff0ef", X"04400513", X"244000ef", X"00048513", X"9c1ff0ef", X"05000513",
        X"234000ef", X"00090513", X"9b1ff0ef", X"00a00513", X"224000ef", X"101007b7", X"00d00713", X"800024b7",
        X"10e78623", X"c0048493", X"0004a503", X"c15ff0ef", X"0004a783", X"80001537", X"da850513", X"00178793",
        X"00f4a023", X"168000ef", X"0004a783", X"0017f793", X"10079a63", X"000054b7", X"5aa48493", X"00000793",
        X"000106b7", X"00179713", X"00f4c633", X"00e68733", X"00c71023", X"00178793", X"fed796e3", X"80001537",
        X"db050513", X"128000ef", X"00000913", X"00010a37", X"01300b13", X"80001cb7", X"80001bb7", X"80001c37",
        X"00141793", X"00fa07b3", X"0084c9b3", X"0007da83", X"01099993", X"0109d993", X"03598a63", X"032b4663",
        X"01091513", X"db8c8593", X"01055513", X"c19ff0ef", X"dbcb8593", X"00098513", X"c0dff0ef", X"d4cc0593",
        X"000a8513", X"c01ff0ef", X"00190913", X"00140413", X"fb4418e3", X"06090e63", X"80001537", X"dc450513",
        X"0ac000ef", X"00090513", X"b39ff0ef", X"00a00513", X"124000ef", X"00042503", X"b29ff0ef", X"00442503",
        X"b21ff0ef", X"00842503", X"b19ff0ef", X"0b812403", X"0bc12083", X"0b412483", X"0b012903", X"0ac12983",
        X"0a812a03", X"0a412a83", X"0a012b03", X"09c12b83", X"09812c03", X"09412c83", X"00a00513", X"0c010113",
        X"0d40006f", X"000104b7", X"fff48493", X"ef1ff06f", X"0b812403", X"0bc12083", X"0b412483", X"0b012903",
        X"0ac12983", X"0a812a03", X"0a412a83", X"0a012b03", X"09c12b83", X"09812c03", X"09412c83", X"80001537",
        X"dd050513", X"0c010113", X"0040006f", X"ff010113", X"00812423", X"00912223", X"00112623", X"00050493",
        X"00000413", X"008487b3", X"0007c503", X"00140413", X"02051663", X"00d00513", X"05c000ef", X"00a00513",
        X"054000ef", X"00c12083", X"00040513", X"00812403", X"00412483", X"01010113", X"00008067", X"038000ef",
        X"fc5ff06f", X"10000737", X"00c74683", X"00d74783", X"00e74503", X"00f74703", X"01869693", X"01079793",
        X"00d7e7b3", X"00e7e7b3", X"00851513", X"00f56533", X"00008067", X"800027b7", X"c047a783", X"ff010113",
        X"00812423", X"00112623", X"00050413", X"00078463", X"000780e7", X"10000737", X"01274783", X"0107f793",
        X"fe079ce3", X"0ff47413", X"00870823", X"00c12083", X"00812403", X"01010113", X"00008067", X"101007b7",
        X"02050063", X"00100713", X"00e785a3", X"101007b7", X"00100713", X"00e78523", X"00078523", X"00008067",
        X"000785a3", X"fe9ff06f", X"ff010113", X"00812423", X"00912223", X"01212023", X"00112623", X"00050493",
        X"00058413", X"02100913", X"00100513", X"fff90913", X"fadff0ef", X"fe091ae3", X"00000513", X"fa1ff0ef",
        X"00100513", X"f99ff0ef", X"00000513", X"f91ff0ef", X"00100513", X"f89ff0ef", X"00000513", X"f81ff0ef",
        X"00000513", X"f79ff0ef", X"00000513", X"f71ff0ef", X"00000513", X"f69ff0ef", X"00000513", X"f61ff0ef",
        X"00500913", X"0104f513", X"fff90913", X"00149493", X"f4dff0ef", X"0ff4f493", X"fe0916e3", X"00100513",
        X"f3dff0ef", X"00000513", X"f35ff0ef", X"01000493", X"ffff8937", X"01247533", X"00141413", X"01041413",
        X"fff48493", X"f19ff0ef", X"01045413", X"fe0494e3", X"00812403", X"00c12083", X"00412483", X"00012903",
        X"00100513", X"01010113", X"ef5ff06f", X"6c6c6548", X"6f77206f", X"2c646c72", X"34365520", X"2149492d",
        X"00000000", X"6967614d", X"000a2163", X"6c707061", X"74616369", X"0a6e6f69", X"00000000", X"6e6e7552",
        X"0a676e69", X"00000000", X"6b636f4c", X"0000000a", X"74706d45", X"77203b79", X"69746961", X"6620676e",
        X"4a20726f", X"20474154", X"67616d69", X"6f742065", X"6f6f6220", X"000a2e74", X"6967614d", X"00203a63",
        X"33323130", X"37363534", X"42413938", X"46454443", X"00000000", X"696c6143", X"74617262", X"206e6f69",
        X"6c696166", X"00006465", X"74697257", X"002e2e65", X"64616552", X"00002e2e", X"0000003a", X"203d2120",
        X"00000000", X"204d4152", X"6f727265", X"000a2e72", X"204d4152", X"21214b4f", X"0000000d", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
        X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000"

    );
end package;
