-- nios.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios is
	port (
		clk50_clk                : in    std_logic                     := '0';             --     clk50.clk
		io_ack                   : in    std_logic                     := '0';             --        io.ack
		io_rdata                 : in    std_logic_vector(7 downto 0)  := (others => '0'); --          .rdata
		io_read                  : out   std_logic;                                        --          .read
		io_wdata                 : out   std_logic_vector(7 downto 0);                     --          .wdata
		io_write                 : out   std_logic;                                        --          .write
		io_address               : out   std_logic_vector(19 downto 0);                    --          .address
		io_irq                   : in    std_logic                     := '0';             --          .irq
		mem32_address            : in    std_logic_vector(25 downto 0) := (others => '0'); --     mem32.address
		mem32_direction          : in    std_logic                     := '0';             --          .direction
		mem32_byte_en            : in    std_logic_vector(3 downto 0)  := (others => '0'); --          .byte_en
		mem32_wdata              : in    std_logic_vector(31 downto 0) := (others => '0'); --          .wdata
		mem32_request            : in    std_logic                     := '0';             --          .request
		mem32_tag                : in    std_logic_vector(7 downto 0)  := (others => '0'); --          .tag
		mem32_dack_tag           : out   std_logic_vector(7 downto 0);                     --          .dack_tag
		mem32_rdata              : out   std_logic_vector(31 downto 0);                    --          .rdata
		mem32_rack               : out   std_logic;                                        --          .rack
		mem32_rack_tag           : out   std_logic_vector(7 downto 0);                     --          .rack_tag
		memory_mem_a             : out   std_logic_vector(13 downto 0);                    --    memory.mem_a
		memory_mem_ba            : out   std_logic_vector(1 downto 0);                     --          .mem_ba
		memory_mem_ck            : out   std_logic_vector(0 downto 0);                     --          .mem_ck
		memory_mem_ck_n          : out   std_logic_vector(0 downto 0);                     --          .mem_ck_n
		memory_mem_cke           : out   std_logic_vector(0 downto 0);                     --          .mem_cke
		memory_mem_cs_n          : out   std_logic_vector(0 downto 0);                     --          .mem_cs_n
		memory_mem_dm            : out   std_logic_vector(0 downto 0);                     --          .mem_dm
		memory_mem_ras_n         : out   std_logic_vector(0 downto 0);                     --          .mem_ras_n
		memory_mem_cas_n         : out   std_logic_vector(0 downto 0);                     --          .mem_cas_n
		memory_mem_we_n          : out   std_logic_vector(0 downto 0);                     --          .mem_we_n
		memory_mem_dq            : inout std_logic_vector(7 downto 0)  := (others => '0'); --          .mem_dq
		memory_mem_dqs           : inout std_logic_vector(0 downto 0)  := (others => '0'); --          .mem_dqs
		memory_mem_dqs_n         : inout std_logic_vector(0 downto 0)  := (others => '0'); --          .mem_dqs_n
		memory_mem_odt           : out   std_logic_vector(0 downto 0);                     --          .mem_odt
		oct_rzqin                : in    std_logic                     := '0';             --       oct.rzqin
		pio_in_port              : in    std_logic_vector(31 downto 0) := (others => '0'); --       pio.in_port
		pio_out_port             : out   std_logic_vector(31 downto 0);                    --          .out_port
		reset_reset_n            : in    std_logic                     := '0';             --     reset.reset_n
		status_local_init_done   : out   std_logic;                                        --    status.local_init_done
		status_local_cal_success : out   std_logic;                                        --          .local_cal_success
		status_local_cal_fail    : out   std_logic;                                        --          .local_cal_fail
		sys_clock_clk            : out   std_logic;                                        -- sys_clock.clk
		sys_reset_reset_n        : out   std_logic                                         -- sys_reset.reset_n
	);
end entity nios;

architecture rtl of nios is
	component avalon_to_io_bridge is
		port (
			reset             : in  std_logic                     := 'X';             -- reset
			avs_read          : in  std_logic                     := 'X';             -- read
			avs_write         : in  std_logic                     := 'X';             -- write
			avs_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			avs_writedata     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			avs_ready         : out std_logic;                                        -- waitrequest_n
			avs_readdata      : out std_logic_vector(7 downto 0);                     -- readdata
			avs_readdatavalid : out std_logic;                                        -- readdatavalid
			clock             : in  std_logic                     := 'X';             -- clk
			io_ack            : in  std_logic                     := 'X';             -- ack
			io_rdata          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rdata
			io_read           : out std_logic;                                        -- read
			io_wdata          : out std_logic_vector(7 downto 0);                     -- wdata
			io_write          : out std_logic;                                        -- write
			io_address        : out std_logic_vector(19 downto 0);                    -- address
			io_irq            : in  std_logic                     := 'X';             -- irq
			avs_irq           : out std_logic                                         -- irq
		);
	end component avalon_to_io_bridge;

	component mem32_to_avalon_bridge is
		port (
			reset              : in  std_logic                     := 'X';             -- reset
			clock              : in  std_logic                     := 'X';             -- clk
			memreq_address     : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			memreq_read_writen : in  std_logic                     := 'X';             -- direction
			memreq_byte_en     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byte_en
			memreq_data        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			memreq_request     : in  std_logic                     := 'X';             -- request
			memreq_tag         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- tag
			memresp_dack_tag   : out std_logic_vector(7 downto 0);                     -- dack_tag
			memresp_data       : out std_logic_vector(31 downto 0);                    -- rdata
			memresp_rack       : out std_logic;                                        -- rack
			memresp_rack_tag   : out std_logic_vector(7 downto 0);                     -- rack_tag
			avm_read           : out std_logic;                                        -- read
			avm_write          : out std_logic;                                        -- write
			avm_address        : out std_logic_vector(25 downto 0);                    -- address
			avm_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			avm_byte_enable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_ready          : in  std_logic                     := 'X';             -- waitrequest_n
			avm_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_readdatavalid  : in  std_logic                     := 'X'              -- readdatavalid
		);
	end component mem32_to_avalon_bridge;

	component nios_mem_if_ddr2_emif_0 is
		port (
			pll_ref_clk        : in    std_logic                     := 'X';             -- clk
			global_reset_n     : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n       : in    std_logic                     := 'X';             -- reset_n
			afi_clk            : out   std_logic;                                        -- clk
			afi_half_clk       : out   std_logic;                                        -- clk
			afi_reset_n        : out   std_logic;                                        -- reset_n
			afi_reset_export_n : out   std_logic;                                        -- reset_n
			mem_a              : out   std_logic_vector(13 downto 0);                    -- mem_a
			mem_ba             : out   std_logic_vector(1 downto 0);                     -- mem_ba
			mem_ck             : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n           : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke            : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n           : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm             : out   std_logic_vector(0 downto 0);                     -- mem_dm
			mem_ras_n          : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			mem_cas_n          : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			mem_we_n           : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			mem_dq             : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs            : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n          : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt            : out   std_logic_vector(0 downto 0);                     -- mem_odt
			avl_ready          : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin     : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr           : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			avl_rdata_valid    : out   std_logic;                                        -- readdatavalid
			avl_rdata          : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata          : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be             : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req       : in    std_logic                     := 'X';             -- read
			avl_write_req      : in    std_logic                     := 'X';             -- write
			avl_size           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			local_init_done    : out   std_logic;                                        -- local_init_done
			local_cal_success  : out   std_logic;                                        -- local_cal_success
			local_cal_fail     : out   std_logic;                                        -- local_cal_fail
			oct_rzqin          : in    std_logic                     := 'X'              -- rzqin
		);
	end component nios_mem_if_ddr2_emif_0;

	component nios_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(28 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_nios2_gen2_0;

	component nios_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			out_port   : out std_logic_vector(31 downto 0);                    -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_pio_0;

	component nios_mm_interconnect_0 is
		port (
			mem_if_ddr2_emif_0_afi_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			mem32_to_avalon_0_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			mem_if_ddr2_emif_0_avl_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mem_if_ddr2_emif_0_soft_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			mem32_to_avalon_0_avalon_master_address                             : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			mem32_to_avalon_0_avalon_master_waitrequest                         : out std_logic;                                        -- waitrequest
			mem32_to_avalon_0_avalon_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mem32_to_avalon_0_avalon_master_read                                : in  std_logic                     := 'X';             -- read
			mem32_to_avalon_0_avalon_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			mem32_to_avalon_0_avalon_master_readdatavalid                       : out std_logic;                                        -- readdatavalid
			mem32_to_avalon_0_avalon_master_write                               : in  std_logic                     := 'X';             -- write
			mem32_to_avalon_0_avalon_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_address                                    : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                                : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                       : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                                      : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                             : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                         : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                                : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			io_bridge_0_avalon_slave_0_address                                  : out std_logic_vector(19 downto 0);                    -- address
			io_bridge_0_avalon_slave_0_write                                    : out std_logic;                                        -- write
			io_bridge_0_avalon_slave_0_read                                     : out std_logic;                                        -- read
			io_bridge_0_avalon_slave_0_readdata                                 : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			io_bridge_0_avalon_slave_0_writedata                                : out std_logic_vector(7 downto 0);                     -- writedata
			io_bridge_0_avalon_slave_0_readdatavalid                            : in  std_logic                     := 'X';             -- readdatavalid
			io_bridge_0_avalon_slave_0_waitrequest                              : in  std_logic                     := 'X';             -- waitrequest
			mem_if_ddr2_emif_0_avl_address                                      : out std_logic_vector(23 downto 0);                    -- address
			mem_if_ddr2_emif_0_avl_write                                        : out std_logic;                                        -- write
			mem_if_ddr2_emif_0_avl_read                                         : out std_logic;                                        -- read
			mem_if_ddr2_emif_0_avl_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mem_if_ddr2_emif_0_avl_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			mem_if_ddr2_emif_0_avl_beginbursttransfer                           : out std_logic;                                        -- beginbursttransfer
			mem_if_ddr2_emif_0_avl_burstcount                                   : out std_logic_vector(2 downto 0);                     -- burstcount
			mem_if_ddr2_emif_0_avl_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			mem_if_ddr2_emif_0_avl_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			mem_if_ddr2_emif_0_avl_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address                                : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                                  : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                                   : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                            : out std_logic;                                        -- debugaccess
			pio_0_s1_address                                                    : out std_logic_vector(2 downto 0);                     -- address
			pio_0_s1_write                                                      : out std_logic;                                        -- write
			pio_0_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                                 : out std_logic                                         -- chipselect
		);
	end component nios_mm_interconnect_0;

	component nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_irq_mapper;

	component nios_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller;

	component nios_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller_001;

	component nios_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller_002;

	signal mem_if_ddr2_emif_0_afi_clk_clk                                : std_logic;                     -- mem_if_ddr2_emif_0:afi_clk -> [sys_clock_clk, io_bridge_0:clock, irq_mapper:clk, mem32_to_avalon_0:clock, mm_interconnect_0:mem_if_ddr2_emif_0_afi_clk_clk, nios2_gen2_0:clk, pio_0:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	signal mm_interconnect_0_mem32_to_avalon_0_avalon_master_waitrequest : std_logic;                     -- mm_interconnect_0:mem32_to_avalon_0_avalon_master_waitrequest -> mm_interconnect_0_mem32_to_avalon_0_avalon_master_waitrequest:in
	signal mem32_to_avalon_0_avalon_master_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:mem32_to_avalon_0_avalon_master_readdata -> mem32_to_avalon_0:avm_readdata
	signal mem32_to_avalon_0_avalon_master_read                          : std_logic;                     -- mem32_to_avalon_0:avm_read -> mm_interconnect_0:mem32_to_avalon_0_avalon_master_read
	signal mem32_to_avalon_0_avalon_master_address                       : std_logic_vector(25 downto 0); -- mem32_to_avalon_0:avm_address -> mm_interconnect_0:mem32_to_avalon_0_avalon_master_address
	signal mem32_to_avalon_0_avalon_master_byteenable                    : std_logic_vector(3 downto 0);  -- mem32_to_avalon_0:avm_byte_enable -> mm_interconnect_0:mem32_to_avalon_0_avalon_master_byteenable
	signal mem32_to_avalon_0_avalon_master_readdatavalid                 : std_logic;                     -- mm_interconnect_0:mem32_to_avalon_0_avalon_master_readdatavalid -> mem32_to_avalon_0:avm_readdatavalid
	signal mem32_to_avalon_0_avalon_master_write                         : std_logic;                     -- mem32_to_avalon_0:avm_write -> mm_interconnect_0:mem32_to_avalon_0_avalon_master_write
	signal mem32_to_avalon_0_avalon_master_writedata                     : std_logic_vector(31 downto 0); -- mem32_to_avalon_0:avm_writedata -> mm_interconnect_0:mem32_to_avalon_0_avalon_master_writedata
	signal nios2_gen2_0_data_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                          : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                              : std_logic_vector(28 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                           : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                 : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                            : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                       : std_logic_vector(28 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                          : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_beginbursttransfer   : std_logic;                     -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_beginbursttransfer -> mem_if_ddr2_emif_0:avl_burstbegin
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdata             : std_logic_vector(31 downto 0); -- mem_if_ddr2_emif_0:avl_rdata -> mm_interconnect_0:mem_if_ddr2_emif_0_avl_readdata
	signal mem_if_ddr2_emif_0_avl_waitrequest                            : std_logic;                     -- mem_if_ddr2_emif_0:avl_ready -> mem_if_ddr2_emif_0_avl_waitrequest:in
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_address              : std_logic_vector(23 downto 0); -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_address -> mem_if_ddr2_emif_0:avl_addr
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_read                 : std_logic;                     -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_read -> mem_if_ddr2_emif_0:avl_read_req
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_byteenable -> mem_if_ddr2_emif_0:avl_be
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdatavalid        : std_logic;                     -- mem_if_ddr2_emif_0:avl_rdata_valid -> mm_interconnect_0:mem_if_ddr2_emif_0_avl_readdatavalid
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_write                : std_logic;                     -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_write -> mem_if_ddr2_emif_0:avl_write_req
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_writedata -> mem_if_ddr2_emif_0:avl_wdata
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_burstcount           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:mem_if_ddr2_emif_0_avl_burstcount -> mem_if_ddr2_emif_0:avl_size
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata       : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest    : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read           : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata         : std_logic_vector(7 downto 0);  -- io_bridge_0:avs_readdata -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdata
	signal io_bridge_0_avalon_slave_0_waitrequest                        : std_logic;                     -- io_bridge_0:avs_ready -> io_bridge_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_address          : std_logic_vector(19 downto 0); -- mm_interconnect_0:io_bridge_0_avalon_slave_0_address -> io_bridge_0:avs_address
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_read             : std_logic;                     -- mm_interconnect_0:io_bridge_0_avalon_slave_0_read -> io_bridge_0:avs_read
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid    : std_logic;                     -- io_bridge_0:avs_readdatavalid -> mm_interconnect_0:io_bridge_0_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:io_bridge_0_avalon_slave_0_write -> io_bridge_0:avs_write
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:io_bridge_0_avalon_slave_0_writedata -> io_bridge_0:avs_writedata
	signal mm_interconnect_0_pio_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                           : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                              : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- io_bridge_0:avs_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- pio_0:irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [io_bridge_0:reset, mem32_to_avalon_0:reset, mm_interconnect_0:mem32_to_avalon_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal mem_if_ddr2_emif_0_afi_reset_reset                            : std_logic;                     -- mem_if_ddr2_emif_0:afi_reset_n -> mem_if_ddr2_emif_0_afi_reset_reset:in
	signal nios2_gen2_0_debug_reset_request_reset                        : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                     -- rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:mem_if_ddr2_emif_0_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr2_emif_0_soft_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller_002:reset_in0
	signal mem32_to_avalon_0_avalon_master_inv                           : std_logic;                     -- mm_interconnect_0_mem32_to_avalon_0_avalon_master_waitrequest:inv -> mem32_to_avalon_0:avm_ready
	signal mm_interconnect_0_mem_if_ddr2_emif_0_avl_inv                  : std_logic;                     -- mem_if_ddr2_emif_0_avl_waitrequest:inv -> mm_interconnect_0:mem_if_ddr2_emif_0_avl_waitrequest
	signal mm_interconnect_0_io_bridge_0_avalon_slave_0_inv              : std_logic;                     -- io_bridge_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:io_bridge_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [sys_reset_reset_n, pio_0:reset_n]
	signal mem_if_ddr2_emif_0_afi_reset_reset_ports_inv                  : std_logic;                     -- mem_if_ddr2_emif_0_afi_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> nios2_gen2_0:reset_n

begin

	io_bridge_0 : component avalon_to_io_bridge
		port map (
			reset             => rst_controller_reset_out_reset,                             --          reset.reset
			avs_read          => mm_interconnect_0_io_bridge_0_avalon_slave_0_read,          -- avalon_slave_0.read
			avs_write         => mm_interconnect_0_io_bridge_0_avalon_slave_0_write,         --               .write
			avs_address       => mm_interconnect_0_io_bridge_0_avalon_slave_0_address,       --               .address
			avs_writedata     => mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata,     --               .writedata
			avs_ready         => io_bridge_0_avalon_slave_0_waitrequest,                     --               .waitrequest_n
			avs_readdata      => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata,      --               .readdata
			avs_readdatavalid => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid, --               .readdatavalid
			clock             => mem_if_ddr2_emif_0_afi_clk_clk,                             --          clock.clk
			io_ack            => io_ack,                                                     --             io.ack
			io_rdata          => io_rdata,                                                   --               .rdata
			io_read           => io_read,                                                    --               .read
			io_wdata          => io_wdata,                                                   --               .wdata
			io_write          => io_write,                                                   --               .write
			io_address        => io_address,                                                 --               .address
			io_irq            => io_irq,                                                     --               .irq
			avs_irq           => irq_mapper_receiver0_irq                                    --            irq.irq
		);

	mem32_to_avalon_0 : component mem32_to_avalon_bridge
		port map (
			reset              => rst_controller_reset_out_reset,                --         reset.reset
			clock              => mem_if_ddr2_emif_0_afi_clk_clk,                --         clock.clk
			memreq_address     => mem32_address,                                 --   mem32_slave.address
			memreq_read_writen => mem32_direction,                               --              .direction
			memreq_byte_en     => mem32_byte_en,                                 --              .byte_en
			memreq_data        => mem32_wdata,                                   --              .wdata
			memreq_request     => mem32_request,                                 --              .request
			memreq_tag         => mem32_tag,                                     --              .tag
			memresp_dack_tag   => mem32_dack_tag,                                --              .dack_tag
			memresp_data       => mem32_rdata,                                   --              .rdata
			memresp_rack       => mem32_rack,                                    --              .rack
			memresp_rack_tag   => mem32_rack_tag,                                --              .rack_tag
			avm_read           => mem32_to_avalon_0_avalon_master_read,          -- avalon_master.read
			avm_write          => mem32_to_avalon_0_avalon_master_write,         --              .write
			avm_address        => mem32_to_avalon_0_avalon_master_address,       --              .address
			avm_writedata      => mem32_to_avalon_0_avalon_master_writedata,     --              .writedata
			avm_byte_enable    => mem32_to_avalon_0_avalon_master_byteenable,    --              .byteenable
			avm_ready          => mem32_to_avalon_0_avalon_master_inv,           --              .waitrequest_n
			avm_readdata       => mem32_to_avalon_0_avalon_master_readdata,      --              .readdata
			avm_readdatavalid  => mem32_to_avalon_0_avalon_master_readdatavalid  --              .readdatavalid
		);

	mem_if_ddr2_emif_0 : component nios_mem_if_ddr2_emif_0
		port map (
			pll_ref_clk        => clk50_clk,                                                   --      pll_ref_clk.clk
			global_reset_n     => reset_reset_n,                                               --     global_reset.reset_n
			soft_reset_n       => reset_reset_n,                                               --       soft_reset.reset_n
			afi_clk            => mem_if_ddr2_emif_0_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk       => open,                                                        --     afi_half_clk.clk
			afi_reset_n        => mem_if_ddr2_emif_0_afi_reset_reset,                          --        afi_reset.reset_n
			afi_reset_export_n => open,                                                        -- afi_reset_export.reset_n
			mem_a              => memory_mem_a,                                                --           memory.mem_a
			mem_ba             => memory_mem_ba,                                               --                 .mem_ba
			mem_ck             => memory_mem_ck,                                               --                 .mem_ck
			mem_ck_n           => memory_mem_ck_n,                                             --                 .mem_ck_n
			mem_cke            => memory_mem_cke,                                              --                 .mem_cke
			mem_cs_n           => memory_mem_cs_n,                                             --                 .mem_cs_n
			mem_dm             => memory_mem_dm,                                               --                 .mem_dm
			mem_ras_n          => memory_mem_ras_n,                                            --                 .mem_ras_n
			mem_cas_n          => memory_mem_cas_n,                                            --                 .mem_cas_n
			mem_we_n           => memory_mem_we_n,                                             --                 .mem_we_n
			mem_dq             => memory_mem_dq,                                               --                 .mem_dq
			mem_dqs            => memory_mem_dqs,                                              --                 .mem_dqs
			mem_dqs_n          => memory_mem_dqs_n,                                            --                 .mem_dqs_n
			mem_odt            => memory_mem_odt,                                              --                 .mem_odt
			avl_ready          => mem_if_ddr2_emif_0_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin     => mm_interconnect_0_mem_if_ddr2_emif_0_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr           => mm_interconnect_0_mem_if_ddr2_emif_0_avl_address,            --                 .address
			avl_rdata_valid    => mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata          => mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdata,           --                 .readdata
			avl_wdata          => mm_interconnect_0_mem_if_ddr2_emif_0_avl_writedata,          --                 .writedata
			avl_be             => mm_interconnect_0_mem_if_ddr2_emif_0_avl_byteenable,         --                 .byteenable
			avl_read_req       => mm_interconnect_0_mem_if_ddr2_emif_0_avl_read,               --                 .read
			avl_write_req      => mm_interconnect_0_mem_if_ddr2_emif_0_avl_write,              --                 .write
			avl_size           => mm_interconnect_0_mem_if_ddr2_emif_0_avl_burstcount,         --                 .burstcount
			local_init_done    => status_local_init_done,                                      --           status.local_init_done
			local_cal_success  => status_local_cal_success,                                    --                 .local_cal_success
			local_cal_fail     => status_local_cal_fail,                                       --                 .local_cal_fail
			oct_rzqin          => oct_rzqin                                                    --              oct.rzqin
		);

	nios2_gen2_0 : component nios_nios2_gen2_0
		port map (
			clk                                 => mem_if_ddr2_emif_0_afi_clk_clk,                             --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	pio_0 : component nios_pio_0
		port map (
			clk        => mem_if_ddr2_emif_0_afi_clk_clk,             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			in_port    => pio_in_port,                                -- external_connection.export
			out_port   => pio_out_port,                               --                    .export
			irq        => irq_mapper_receiver1_irq                    --                 irq.irq
		);

	mm_interconnect_0 : component nios_mm_interconnect_0
		port map (
			mem_if_ddr2_emif_0_afi_clk_clk                                      => mem_if_ddr2_emif_0_afi_clk_clk,                                --                                    mem_if_ddr2_emif_0_afi_clk.clk
			mem32_to_avalon_0_reset_reset_bridge_in_reset_reset                 => rst_controller_reset_out_reset,                                --                 mem32_to_avalon_0_reset_reset_bridge_in_reset.reset
			mem_if_ddr2_emif_0_avl_translator_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                            -- mem_if_ddr2_emif_0_avl_translator_reset_reset_bridge_in_reset.reset
			mem_if_ddr2_emif_0_soft_reset_reset_bridge_in_reset_reset           => rst_controller_002_reset_out_reset,                            --           mem_if_ddr2_emif_0_soft_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                      => rst_controller_001_reset_out_reset,                            --                      nios2_gen2_0_reset_reset_bridge_in_reset.reset
			mem32_to_avalon_0_avalon_master_address                             => mem32_to_avalon_0_avalon_master_address,                       --                               mem32_to_avalon_0_avalon_master.address
			mem32_to_avalon_0_avalon_master_waitrequest                         => mm_interconnect_0_mem32_to_avalon_0_avalon_master_waitrequest, --                                                              .waitrequest
			mem32_to_avalon_0_avalon_master_byteenable                          => mem32_to_avalon_0_avalon_master_byteenable,                    --                                                              .byteenable
			mem32_to_avalon_0_avalon_master_read                                => mem32_to_avalon_0_avalon_master_read,                          --                                                              .read
			mem32_to_avalon_0_avalon_master_readdata                            => mem32_to_avalon_0_avalon_master_readdata,                      --                                                              .readdata
			mem32_to_avalon_0_avalon_master_readdatavalid                       => mem32_to_avalon_0_avalon_master_readdatavalid,                 --                                                              .readdatavalid
			mem32_to_avalon_0_avalon_master_write                               => mem32_to_avalon_0_avalon_master_write,                         --                                                              .write
			mem32_to_avalon_0_avalon_master_writedata                           => mem32_to_avalon_0_avalon_master_writedata,                     --                                                              .writedata
			nios2_gen2_0_data_master_address                                    => nios2_gen2_0_data_master_address,                              --                                      nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                                => nios2_gen2_0_data_master_waitrequest,                          --                                                              .waitrequest
			nios2_gen2_0_data_master_byteenable                                 => nios2_gen2_0_data_master_byteenable,                           --                                                              .byteenable
			nios2_gen2_0_data_master_read                                       => nios2_gen2_0_data_master_read,                                 --                                                              .read
			nios2_gen2_0_data_master_readdata                                   => nios2_gen2_0_data_master_readdata,                             --                                                              .readdata
			nios2_gen2_0_data_master_write                                      => nios2_gen2_0_data_master_write,                                --                                                              .write
			nios2_gen2_0_data_master_writedata                                  => nios2_gen2_0_data_master_writedata,                            --                                                              .writedata
			nios2_gen2_0_data_master_debugaccess                                => nios2_gen2_0_data_master_debugaccess,                          --                                                              .debugaccess
			nios2_gen2_0_instruction_master_address                             => nios2_gen2_0_instruction_master_address,                       --                               nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                         => nios2_gen2_0_instruction_master_waitrequest,                   --                                                              .waitrequest
			nios2_gen2_0_instruction_master_read                                => nios2_gen2_0_instruction_master_read,                          --                                                              .read
			nios2_gen2_0_instruction_master_readdata                            => nios2_gen2_0_instruction_master_readdata,                      --                                                              .readdata
			io_bridge_0_avalon_slave_0_address                                  => mm_interconnect_0_io_bridge_0_avalon_slave_0_address,          --                                    io_bridge_0_avalon_slave_0.address
			io_bridge_0_avalon_slave_0_write                                    => mm_interconnect_0_io_bridge_0_avalon_slave_0_write,            --                                                              .write
			io_bridge_0_avalon_slave_0_read                                     => mm_interconnect_0_io_bridge_0_avalon_slave_0_read,             --                                                              .read
			io_bridge_0_avalon_slave_0_readdata                                 => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdata,         --                                                              .readdata
			io_bridge_0_avalon_slave_0_writedata                                => mm_interconnect_0_io_bridge_0_avalon_slave_0_writedata,        --                                                              .writedata
			io_bridge_0_avalon_slave_0_readdatavalid                            => mm_interconnect_0_io_bridge_0_avalon_slave_0_readdatavalid,    --                                                              .readdatavalid
			io_bridge_0_avalon_slave_0_waitrequest                              => mm_interconnect_0_io_bridge_0_avalon_slave_0_inv,              --                                                              .waitrequest
			mem_if_ddr2_emif_0_avl_address                                      => mm_interconnect_0_mem_if_ddr2_emif_0_avl_address,              --                                        mem_if_ddr2_emif_0_avl.address
			mem_if_ddr2_emif_0_avl_write                                        => mm_interconnect_0_mem_if_ddr2_emif_0_avl_write,                --                                                              .write
			mem_if_ddr2_emif_0_avl_read                                         => mm_interconnect_0_mem_if_ddr2_emif_0_avl_read,                 --                                                              .read
			mem_if_ddr2_emif_0_avl_readdata                                     => mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdata,             --                                                              .readdata
			mem_if_ddr2_emif_0_avl_writedata                                    => mm_interconnect_0_mem_if_ddr2_emif_0_avl_writedata,            --                                                              .writedata
			mem_if_ddr2_emif_0_avl_beginbursttransfer                           => mm_interconnect_0_mem_if_ddr2_emif_0_avl_beginbursttransfer,   --                                                              .beginbursttransfer
			mem_if_ddr2_emif_0_avl_burstcount                                   => mm_interconnect_0_mem_if_ddr2_emif_0_avl_burstcount,           --                                                              .burstcount
			mem_if_ddr2_emif_0_avl_byteenable                                   => mm_interconnect_0_mem_if_ddr2_emif_0_avl_byteenable,           --                                                              .byteenable
			mem_if_ddr2_emif_0_avl_readdatavalid                                => mm_interconnect_0_mem_if_ddr2_emif_0_avl_readdatavalid,        --                                                              .readdatavalid
			mem_if_ddr2_emif_0_avl_waitrequest                                  => mm_interconnect_0_mem_if_ddr2_emif_0_avl_inv,                  --                                                              .waitrequest
			nios2_gen2_0_debug_mem_slave_address                                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,        --                                  nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,          --                                                              .write
			nios2_gen2_0_debug_mem_slave_read                                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,           --                                                              .read
			nios2_gen2_0_debug_mem_slave_readdata                               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,       --                                                              .readdata
			nios2_gen2_0_debug_mem_slave_writedata                              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,      --                                                              .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,     --                                                              .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,    --                                                              .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,    --                                                              .debugaccess
			pio_0_s1_address                                                    => mm_interconnect_0_pio_0_s1_address,                            --                                                      pio_0_s1.address
			pio_0_s1_write                                                      => mm_interconnect_0_pio_0_s1_write,                              --                                                              .write
			pio_0_s1_readdata                                                   => mm_interconnect_0_pio_0_s1_readdata,                           --                                                              .readdata
			pio_0_s1_writedata                                                  => mm_interconnect_0_pio_0_s1_writedata,                          --                                                              .writedata
			pio_0_s1_chipselect                                                 => mm_interconnect_0_pio_0_s1_chipselect                          --                                                              .chipselect
		);

	irq_mapper : component nios_irq_mapper
		port map (
			clk           => mem_if_ddr2_emif_0_afi_clk_clk,     --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	rst_controller : component nios_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => mem_if_ddr2_emif_0_afi_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset,       -- reset_in1.reset
			clk            => mem_if_ddr2_emif_0_afi_clk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,               -- reset_out.reset
			reset_req      => open,                                         -- (terminated)
			reset_req_in0  => '0',                                          -- (terminated)
			reset_req_in1  => '0',                                          -- (terminated)
			reset_in2      => '0',                                          -- (terminated)
			reset_req_in2  => '0',                                          -- (terminated)
			reset_in3      => '0',                                          -- (terminated)
			reset_req_in3  => '0',                                          -- (terminated)
			reset_in4      => '0',                                          -- (terminated)
			reset_req_in4  => '0',                                          -- (terminated)
			reset_in5      => '0',                                          -- (terminated)
			reset_req_in5  => '0',                                          -- (terminated)
			reset_in6      => '0',                                          -- (terminated)
			reset_req_in6  => '0',                                          -- (terminated)
			reset_in7      => '0',                                          -- (terminated)
			reset_req_in7  => '0',                                          -- (terminated)
			reset_in8      => '0',                                          -- (terminated)
			reset_req_in8  => '0',                                          -- (terminated)
			reset_in9      => '0',                                          -- (terminated)
			reset_req_in9  => '0',                                          -- (terminated)
			reset_in10     => '0',                                          -- (terminated)
			reset_req_in10 => '0',                                          -- (terminated)
			reset_in11     => '0',                                          -- (terminated)
			reset_req_in11 => '0',                                          -- (terminated)
			reset_in12     => '0',                                          -- (terminated)
			reset_req_in12 => '0',                                          -- (terminated)
			reset_in13     => '0',                                          -- (terminated)
			reset_req_in13 => '0',                                          -- (terminated)
			reset_in14     => '0',                                          -- (terminated)
			reset_req_in14 => '0',                                          -- (terminated)
			reset_in15     => '0',                                          -- (terminated)
			reset_req_in15 => '0'                                           -- (terminated)
		);

	rst_controller_001 : component nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => mem_if_ddr2_emif_0_afi_reset_reset_ports_inv, -- reset_in0.reset
			clk            => mem_if_ddr2_emif_0_afi_clk_clk,               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,           -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,       --          .reset_req
			reset_req_in0  => '0',                                          -- (terminated)
			reset_in1      => '0',                                          -- (terminated)
			reset_req_in1  => '0',                                          -- (terminated)
			reset_in2      => '0',                                          -- (terminated)
			reset_req_in2  => '0',                                          -- (terminated)
			reset_in3      => '0',                                          -- (terminated)
			reset_req_in3  => '0',                                          -- (terminated)
			reset_in4      => '0',                                          -- (terminated)
			reset_req_in4  => '0',                                          -- (terminated)
			reset_in5      => '0',                                          -- (terminated)
			reset_req_in5  => '0',                                          -- (terminated)
			reset_in6      => '0',                                          -- (terminated)
			reset_req_in6  => '0',                                          -- (terminated)
			reset_in7      => '0',                                          -- (terminated)
			reset_req_in7  => '0',                                          -- (terminated)
			reset_in8      => '0',                                          -- (terminated)
			reset_req_in8  => '0',                                          -- (terminated)
			reset_in9      => '0',                                          -- (terminated)
			reset_req_in9  => '0',                                          -- (terminated)
			reset_in10     => '0',                                          -- (terminated)
			reset_req_in10 => '0',                                          -- (terminated)
			reset_in11     => '0',                                          -- (terminated)
			reset_req_in11 => '0',                                          -- (terminated)
			reset_in12     => '0',                                          -- (terminated)
			reset_req_in12 => '0',                                          -- (terminated)
			reset_in13     => '0',                                          -- (terminated)
			reset_req_in13 => '0',                                          -- (terminated)
			reset_in14     => '0',                                          -- (terminated)
			reset_req_in14 => '0',                                          -- (terminated)
			reset_in15     => '0',                                          -- (terminated)
			reset_req_in15 => '0'                                           -- (terminated)
		);

	rst_controller_002 : component nios_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => mem_if_ddr2_emif_0_afi_clk_clk,     --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mem32_to_avalon_0_avalon_master_inv <= not mm_interconnect_0_mem32_to_avalon_0_avalon_master_waitrequest;

	mm_interconnect_0_mem_if_ddr2_emif_0_avl_inv <= not mem_if_ddr2_emif_0_avl_waitrequest;

	mm_interconnect_0_io_bridge_0_avalon_slave_0_inv <= not io_bridge_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	mem_if_ddr2_emif_0_afi_reset_reset_ports_inv <= not mem_if_ddr2_emif_0_afi_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	sys_clock_clk <= mem_if_ddr2_emif_0_afi_clk_clk;

	sys_reset_reset_n <= rst_controller_reset_out_reset_ports_inv;

end architecture rtl; -- of nios
