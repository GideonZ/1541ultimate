
module nios (
	clk_clk,
	reset_reset_n,
	nios2_gen2_0_irq_irq);	

	input		clk_clk;
	input		reset_reset_n;
	input	[31:0]	nios2_gen2_0_irq_irq;
endmodule
